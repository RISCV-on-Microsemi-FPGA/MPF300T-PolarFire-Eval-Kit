`timescale 1 ns/100 ps
// Version: 


module HS_IO_CLK(
       A,
       Y
    )
/* synthesis black_box

pragma attribute HS_IO_CLK ment_tpd0 A->Y+1.384
*/
/* synthesis black_box black_box_pad ="" */
 ;
input  A;
output Y;

endmodule
