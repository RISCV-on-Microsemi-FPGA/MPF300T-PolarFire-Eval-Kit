// Copyright 2009 Actel Corporation. All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// Revision Information:
// SVN Revision Information:
// SVN $Revision: $
module
CAHBtoAPB3O
(
input
wire
HCLK,
input
wire
HRESETN,
input
wire
HSEL,
input
wire
CAHBtoAPB3I,
input
wire
HWRITE,
input
wire
HREADY,
output
reg
[
1
:
0
]
HRESP,
output
reg
HREADYOUT,
input
wire
PREADY,
input
wire
PSLVERR,
input
wire
PENABLE,
output
reg
PWRITE,
output
reg
PSEL,
output
reg
CAHBtoAPB3l,
output
reg
CAHBtoAPB3OI,
output
reg
CAHBtoAPB3II,
output
reg
CAHBtoAPB3lI,
output
reg
CAHBtoAPB3Ol,
output
reg
CAHBtoAPB3Il,
output
reg
CAHBtoAPB3ll
)
;
parameter
SYNC_RESET
=
0
;
localparam
CAHBtoAPB3O0
=
2
'b
00
;
localparam
CAHBtoAPB3I0
=
2
'b
01
;
localparam
CAHBtoAPB3l0
=
3
'b
000
;
localparam
CAHBtoAPB3O1
=
3
'b
001
;
localparam
CAHBtoAPB3I1
=
3
'b
010
;
localparam
CAHBtoAPB3l1
=
3
'b
011
;
localparam
CAHBtoAPB3OOI
=
3
'b
100
;
reg
[
2
:
0
]
CAHBtoAPB3IOI
,
CAHBtoAPB3lOI
;
reg
CAHBtoAPB3OII
;
reg
CAHBtoAPB3III
;
reg
CAHBtoAPB3lII
;
reg
CAHBtoAPB3OlI
;
reg
CAHBtoAPB3IlI
;
reg
CAHBtoAPB3llI
;
reg
CAHBtoAPB3O0I
;
reg
CAHBtoAPB3I0I
;
reg
CAHBtoAPB3l0I
;
wire
CAHBtoAPB3O1I
;
wire
CAHBtoAPB3I1I
;
assign
CAHBtoAPB3O1I
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
HRESETN
;
assign
CAHBtoAPB3I1I
=
(
SYNC_RESET
==
1
)
?
HRESETN
:
1
'b
1
;
always
@
(
*
)
begin
CAHBtoAPB3l
=
1
'b
0
;
CAHBtoAPB3OI
=
1
'b
0
;
CAHBtoAPB3II
=
1
'b
0
;
CAHBtoAPB3lI
=
1
'b
0
;
CAHBtoAPB3OII
=
1
'b
0
;
CAHBtoAPB3Ol
=
1
'b
0
;
CAHBtoAPB3OlI
=
1
'b
0
;
CAHBtoAPB3IlI
=
1
'b
0
;
CAHBtoAPB3Il
=
1
'b
0
;
CAHBtoAPB3ll
=
1
'b
0
;
CAHBtoAPB3llI
=
1
'b
0
;
CAHBtoAPB3O0I
=
1
'b
0
;
CAHBtoAPB3I0I
=
1
'b
1
;
case
(
CAHBtoAPB3IOI
)
CAHBtoAPB3l0
:
begin
if
(
HSEL
&&
HREADY
&&
CAHBtoAPB3I
)
begin
CAHBtoAPB3l
=
1
'b
1
;
if
(
HWRITE
)
begin
CAHBtoAPB3lOI
=
CAHBtoAPB3O1
;
end
else
begin
CAHBtoAPB3Il
=
1
'b
1
;
CAHBtoAPB3llI
=
1
'b
1
;
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lOI
=
CAHBtoAPB3l1
;
end
end
else
begin
CAHBtoAPB3lOI
=
CAHBtoAPB3l0
;
end
end
CAHBtoAPB3O1
:
begin
if
(
HSEL
&&
HREADY
&&
CAHBtoAPB3I
)
begin
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lI
=
1
'b
1
;
CAHBtoAPB3OII
=
1
'b
1
;
CAHBtoAPB3OlI
=
1
'b
1
;
end
CAHBtoAPB3OI
=
1
'b
1
;
CAHBtoAPB3Il
=
1
'b
1
;
CAHBtoAPB3llI
=
1
'b
1
;
CAHBtoAPB3O0I
=
1
'b
1
;
CAHBtoAPB3lOI
=
CAHBtoAPB3I1
;
end
CAHBtoAPB3I1
:
begin
if
(
PENABLE
&&
PREADY
)
begin
CAHBtoAPB3ll
=
1
'b
1
;
if
(
HSEL
&&
HREADY
&&
CAHBtoAPB3I
)
begin
CAHBtoAPB3l
=
1
'b
1
;
if
(
HWRITE
)
begin
CAHBtoAPB3lOI
=
CAHBtoAPB3O1
;
end
else
begin
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lOI
=
CAHBtoAPB3OOI
;
end
end
else
begin
if
(
CAHBtoAPB3lII
)
begin
CAHBtoAPB3Ol
=
1
'b
1
;
CAHBtoAPB3IlI
=
1
'b
1
;
if
(
CAHBtoAPB3III
)
begin
CAHBtoAPB3lOI
=
CAHBtoAPB3O1
;
end
else
begin
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lOI
=
CAHBtoAPB3OOI
;
end
end
else
begin
CAHBtoAPB3lOI
=
CAHBtoAPB3l0
;
end
end
end
else
begin
CAHBtoAPB3llI
=
1
'b
1
;
CAHBtoAPB3O0I
=
1
'b
1
;
if
(
CAHBtoAPB3lII
)
begin
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lOI
=
CAHBtoAPB3I1
;
end
else
begin
if
(
HSEL
&&
HREADY
&&
CAHBtoAPB3I
)
begin
CAHBtoAPB3lI
=
1
'b
1
;
CAHBtoAPB3OII
=
1
'b
1
;
CAHBtoAPB3OlI
=
1
'b
1
;
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lOI
=
CAHBtoAPB3I1
;
end
else
begin
CAHBtoAPB3lOI
=
CAHBtoAPB3I1
;
end
end
end
end
CAHBtoAPB3l1
:
begin
if
(
PENABLE
&&
PREADY
)
begin
CAHBtoAPB3II
=
1
'b
1
;
CAHBtoAPB3ll
=
1
'b
1
;
CAHBtoAPB3lOI
=
CAHBtoAPB3l0
;
end
else
begin
CAHBtoAPB3llI
=
1
'b
1
;
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lOI
=
CAHBtoAPB3l1
;
end
end
CAHBtoAPB3OOI
:
begin
CAHBtoAPB3Il
=
1
'b
1
;
CAHBtoAPB3llI
=
1
'b
1
;
CAHBtoAPB3I0I
=
1
'b
0
;
CAHBtoAPB3lOI
=
CAHBtoAPB3l1
;
end
default
:
begin
CAHBtoAPB3lOI
=
CAHBtoAPB3l0
;
end
endcase
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3IOI
<=
CAHBtoAPB3l0
;
PSEL
<=
1
'b
0
;
PWRITE
<=
1
'b
0
;
end
else
begin
CAHBtoAPB3IOI
<=
CAHBtoAPB3lOI
;
PSEL
<=
CAHBtoAPB3llI
;
PWRITE
<=
CAHBtoAPB3O0I
;
end
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3lII
<=
1
'b
0
;
end
else
begin
if
(
CAHBtoAPB3OlI
)
begin
CAHBtoAPB3lII
<=
1
'b
1
;
end
else
begin
if
(
CAHBtoAPB3IlI
)
begin
CAHBtoAPB3lII
<=
1
'b
0
;
end
end
end
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3III
<=
1
'b
0
;
end
else
begin
if
(
CAHBtoAPB3OII
)
begin
CAHBtoAPB3III
<=
HWRITE
;
end
end
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3l0I
<=
1
'b
0
;
HRESP
<=
CAHBtoAPB3O0
;
HREADYOUT
<=
1
'b
1
;
end
else
begin
case
(
CAHBtoAPB3l0I
)
1
'b
0
:
begin
if
(
PSLVERR
)
begin
CAHBtoAPB3l0I
<=
1
'b
1
;
HRESP
<=
CAHBtoAPB3I0
;
HREADYOUT
<=
1
'b
0
;
end
else
begin
CAHBtoAPB3l0I
<=
1
'b
0
;
HRESP
<=
CAHBtoAPB3O0
;
HREADYOUT
<=
CAHBtoAPB3I0I
;
end
end
1
'b
1
:
begin
CAHBtoAPB3l0I
<=
1
'b
0
;
HRESP
<=
CAHBtoAPB3I0
;
HREADYOUT
<=
1
'b
1
;
end
default
:
begin
CAHBtoAPB3l0I
<=
1
'b
0
;
end
endcase
end
end
endmodule
