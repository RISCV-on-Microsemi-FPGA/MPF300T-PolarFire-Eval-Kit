`timescale 1 ns/100 ps
// Version: 


module HS_IO_CLK(
       A,
       Y
    ) ;
/* synthesis syn_black_box

syn_tpd0 = " A->Y = 1.384"
*/
/* synthesis black_box_pad_pin ="" */
input  A;
output Y;

endmodule
