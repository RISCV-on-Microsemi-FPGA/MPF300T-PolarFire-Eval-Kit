`timescale 1 ns/100 ps
// Version: PolarFire v1.1SP1 12.100.9.11


module lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM(
       W_DATA,
       R_DATA,
       W_ADDR,
       R_ADDR,
       W_EN,
       R_EN,
       CLK,
       WBYTE_EN
    );
input  [39:0] W_DATA;
output [39:0] R_DATA;
input  [17:0] W_ADDR;
input  [17:0] R_ADDR;
input  W_EN;
input  R_EN;
input  CLK;
input  [19:0] WBYTE_EN;

    wire \R_DATA_TEMPR0[0] , \R_DATA_TEMPR1[0] , \R_DATA_TEMPR2[0] , 
        \R_DATA_TEMPR3[0] , \R_DATA_TEMPR4[0] , \R_DATA_TEMPR5[0] , 
        \R_DATA_TEMPR6[0] , \R_DATA_TEMPR7[0] , \R_DATA_TEMPR8[0] , 
        \R_DATA_TEMPR9[0] , \R_DATA_TEMPR10[0] , \R_DATA_TEMPR11[0] , 
        \R_DATA_TEMPR12[0] , \R_DATA_TEMPR13[0] , \R_DATA_TEMPR14[0] , 
        \R_DATA_TEMPR15[0] , \R_DATA_TEMPR16[0] , \R_DATA_TEMPR17[0] , 
        \R_DATA_TEMPR18[0] , \R_DATA_TEMPR19[0] , \R_DATA_TEMPR20[0] , 
        \R_DATA_TEMPR21[0] , \R_DATA_TEMPR22[0] , \R_DATA_TEMPR23[0] , 
        \R_DATA_TEMPR24[0] , \R_DATA_TEMPR25[0] , \R_DATA_TEMPR26[0] , 
        \R_DATA_TEMPR27[0] , \R_DATA_TEMPR28[0] , \R_DATA_TEMPR29[0] , 
        \R_DATA_TEMPR30[0] , \R_DATA_TEMPR31[0] , \R_DATA_TEMPR0[1] , 
        \R_DATA_TEMPR1[1] , \R_DATA_TEMPR2[1] , \R_DATA_TEMPR3[1] , 
        \R_DATA_TEMPR4[1] , \R_DATA_TEMPR5[1] , \R_DATA_TEMPR6[1] , 
        \R_DATA_TEMPR7[1] , \R_DATA_TEMPR8[1] , \R_DATA_TEMPR9[1] , 
        \R_DATA_TEMPR10[1] , \R_DATA_TEMPR11[1] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR13[1] , \R_DATA_TEMPR14[1] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR16[1] , \R_DATA_TEMPR17[1] , \R_DATA_TEMPR18[1] , 
        \R_DATA_TEMPR19[1] , \R_DATA_TEMPR20[1] , \R_DATA_TEMPR21[1] , 
        \R_DATA_TEMPR22[1] , \R_DATA_TEMPR23[1] , \R_DATA_TEMPR24[1] , 
        \R_DATA_TEMPR25[1] , \R_DATA_TEMPR26[1] , \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR28[1] , \R_DATA_TEMPR29[1] , \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR31[1] , \R_DATA_TEMPR0[2] , \R_DATA_TEMPR1[2] , 
        \R_DATA_TEMPR2[2] , \R_DATA_TEMPR3[2] , \R_DATA_TEMPR4[2] , 
        \R_DATA_TEMPR5[2] , \R_DATA_TEMPR6[2] , \R_DATA_TEMPR7[2] , 
        \R_DATA_TEMPR8[2] , \R_DATA_TEMPR9[2] , \R_DATA_TEMPR10[2] , 
        \R_DATA_TEMPR11[2] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR13[2] , 
        \R_DATA_TEMPR14[2] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR16[2] , 
        \R_DATA_TEMPR17[2] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR19[2] , 
        \R_DATA_TEMPR20[2] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR22[2] , 
        \R_DATA_TEMPR23[2] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR25[2] , 
        \R_DATA_TEMPR26[2] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR28[2] , 
        \R_DATA_TEMPR29[2] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR31[2] , 
        \R_DATA_TEMPR0[3] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR2[3] , 
        \R_DATA_TEMPR3[3] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR5[3] , 
        \R_DATA_TEMPR6[3] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR8[3] , 
        \R_DATA_TEMPR9[3] , \R_DATA_TEMPR10[3] , \R_DATA_TEMPR11[3] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR13[3] , \R_DATA_TEMPR14[3] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR16[3] , \R_DATA_TEMPR17[3] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR19[3] , \R_DATA_TEMPR20[3] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR22[3] , \R_DATA_TEMPR23[3] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR25[3] , \R_DATA_TEMPR26[3] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR28[3] , \R_DATA_TEMPR29[3] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR31[3] , \R_DATA_TEMPR0[4] , 
        \R_DATA_TEMPR1[4] , \R_DATA_TEMPR2[4] , \R_DATA_TEMPR3[4] , 
        \R_DATA_TEMPR4[4] , \R_DATA_TEMPR5[4] , \R_DATA_TEMPR6[4] , 
        \R_DATA_TEMPR7[4] , \R_DATA_TEMPR8[4] , \R_DATA_TEMPR9[4] , 
        \R_DATA_TEMPR10[4] , \R_DATA_TEMPR11[4] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR13[4] , \R_DATA_TEMPR14[4] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR16[4] , \R_DATA_TEMPR17[4] , \R_DATA_TEMPR18[4] , 
        \R_DATA_TEMPR19[4] , \R_DATA_TEMPR20[4] , \R_DATA_TEMPR21[4] , 
        \R_DATA_TEMPR22[4] , \R_DATA_TEMPR23[4] , \R_DATA_TEMPR24[4] , 
        \R_DATA_TEMPR25[4] , \R_DATA_TEMPR26[4] , \R_DATA_TEMPR27[4] , 
        \R_DATA_TEMPR28[4] , \R_DATA_TEMPR29[4] , \R_DATA_TEMPR30[4] , 
        \R_DATA_TEMPR31[4] , \R_DATA_TEMPR0[5] , \R_DATA_TEMPR1[5] , 
        \R_DATA_TEMPR2[5] , \R_DATA_TEMPR3[5] , \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR5[5] , \R_DATA_TEMPR6[5] , \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR8[5] , \R_DATA_TEMPR9[5] , \R_DATA_TEMPR10[5] , 
        \R_DATA_TEMPR11[5] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR13[5] , 
        \R_DATA_TEMPR14[5] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR16[5] , 
        \R_DATA_TEMPR17[5] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR19[5] , 
        \R_DATA_TEMPR20[5] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR22[5] , 
        \R_DATA_TEMPR23[5] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR25[5] , 
        \R_DATA_TEMPR26[5] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR28[5] , 
        \R_DATA_TEMPR29[5] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR31[5] , 
        \R_DATA_TEMPR0[6] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR2[6] , 
        \R_DATA_TEMPR3[6] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR5[6] , 
        \R_DATA_TEMPR6[6] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR8[6] , 
        \R_DATA_TEMPR9[6] , \R_DATA_TEMPR10[6] , \R_DATA_TEMPR11[6] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR13[6] , \R_DATA_TEMPR14[6] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR16[6] , \R_DATA_TEMPR17[6] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR19[6] , \R_DATA_TEMPR20[6] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR22[6] , \R_DATA_TEMPR23[6] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR25[6] , \R_DATA_TEMPR26[6] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR28[6] , \R_DATA_TEMPR29[6] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR31[6] , \R_DATA_TEMPR0[7] , 
        \R_DATA_TEMPR1[7] , \R_DATA_TEMPR2[7] , \R_DATA_TEMPR3[7] , 
        \R_DATA_TEMPR4[7] , \R_DATA_TEMPR5[7] , \R_DATA_TEMPR6[7] , 
        \R_DATA_TEMPR7[7] , \R_DATA_TEMPR8[7] , \R_DATA_TEMPR9[7] , 
        \R_DATA_TEMPR10[7] , \R_DATA_TEMPR11[7] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR13[7] , \R_DATA_TEMPR14[7] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR16[7] , \R_DATA_TEMPR17[7] , \R_DATA_TEMPR18[7] , 
        \R_DATA_TEMPR19[7] , \R_DATA_TEMPR20[7] , \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR22[7] , \R_DATA_TEMPR23[7] , \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR25[7] , \R_DATA_TEMPR26[7] , \R_DATA_TEMPR27[7] , 
        \R_DATA_TEMPR28[7] , \R_DATA_TEMPR29[7] , \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR31[7] , \R_DATA_TEMPR0[8] , \R_DATA_TEMPR1[8] , 
        \R_DATA_TEMPR2[8] , \R_DATA_TEMPR3[8] , \R_DATA_TEMPR4[8] , 
        \R_DATA_TEMPR5[8] , \R_DATA_TEMPR6[8] , \R_DATA_TEMPR7[8] , 
        \R_DATA_TEMPR8[8] , \R_DATA_TEMPR9[8] , \R_DATA_TEMPR10[8] , 
        \R_DATA_TEMPR11[8] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR13[8] , 
        \R_DATA_TEMPR14[8] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR16[8] , 
        \R_DATA_TEMPR17[8] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR19[8] , 
        \R_DATA_TEMPR20[8] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR22[8] , 
        \R_DATA_TEMPR23[8] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR25[8] , 
        \R_DATA_TEMPR26[8] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR28[8] , 
        \R_DATA_TEMPR29[8] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR31[8] , 
        \R_DATA_TEMPR0[9] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR2[9] , 
        \R_DATA_TEMPR3[9] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR5[9] , 
        \R_DATA_TEMPR6[9] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR8[9] , 
        \R_DATA_TEMPR9[9] , \R_DATA_TEMPR10[9] , \R_DATA_TEMPR11[9] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR13[9] , \R_DATA_TEMPR14[9] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR16[9] , \R_DATA_TEMPR17[9] , 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR19[9] , \R_DATA_TEMPR20[9] , 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR22[9] , \R_DATA_TEMPR23[9] , 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR25[9] , \R_DATA_TEMPR26[9] , 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR28[9] , \R_DATA_TEMPR29[9] , 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR31[9] , \R_DATA_TEMPR0[10] , 
        \R_DATA_TEMPR1[10] , \R_DATA_TEMPR2[10] , \R_DATA_TEMPR3[10] , 
        \R_DATA_TEMPR4[10] , \R_DATA_TEMPR5[10] , \R_DATA_TEMPR6[10] , 
        \R_DATA_TEMPR7[10] , \R_DATA_TEMPR8[10] , \R_DATA_TEMPR9[10] , 
        \R_DATA_TEMPR10[10] , \R_DATA_TEMPR11[10] , 
        \R_DATA_TEMPR12[10] , \R_DATA_TEMPR13[10] , 
        \R_DATA_TEMPR14[10] , \R_DATA_TEMPR15[10] , 
        \R_DATA_TEMPR16[10] , \R_DATA_TEMPR17[10] , 
        \R_DATA_TEMPR18[10] , \R_DATA_TEMPR19[10] , 
        \R_DATA_TEMPR20[10] , \R_DATA_TEMPR21[10] , 
        \R_DATA_TEMPR22[10] , \R_DATA_TEMPR23[10] , 
        \R_DATA_TEMPR24[10] , \R_DATA_TEMPR25[10] , 
        \R_DATA_TEMPR26[10] , \R_DATA_TEMPR27[10] , 
        \R_DATA_TEMPR28[10] , \R_DATA_TEMPR29[10] , 
        \R_DATA_TEMPR30[10] , \R_DATA_TEMPR31[10] , 
        \R_DATA_TEMPR0[11] , \R_DATA_TEMPR1[11] , \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR3[11] , \R_DATA_TEMPR4[11] , \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR6[11] , \R_DATA_TEMPR7[11] , \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR9[11] , \R_DATA_TEMPR10[11] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR12[11] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR14[11] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR16[11] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR18[11] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR20[11] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR22[11] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR24[11] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR26[11] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR28[11] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR30[11] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR1[12] , 
        \R_DATA_TEMPR2[12] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR4[12] , 
        \R_DATA_TEMPR5[12] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR7[12] , 
        \R_DATA_TEMPR8[12] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR11[12] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR13[12] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR15[12] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR17[12] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR19[12] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR21[12] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR23[12] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR25[12] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR27[12] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR29[12] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR31[12] , \R_DATA_TEMPR0[13] , \R_DATA_TEMPR1[13] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR3[13] , \R_DATA_TEMPR4[13] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR6[13] , \R_DATA_TEMPR7[13] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR9[13] , \R_DATA_TEMPR10[13] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR12[13] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR14[13] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR16[13] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR18[13] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR20[13] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR22[13] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR24[13] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR26[13] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR28[13] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR30[13] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR0[14] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR2[14] , \R_DATA_TEMPR3[14] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR5[14] , \R_DATA_TEMPR6[14] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR8[14] , \R_DATA_TEMPR9[14] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR11[14] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR13[14] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR15[14] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR17[14] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR19[14] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR21[14] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR23[14] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR25[14] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR27[14] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR29[14] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR31[14] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR1[15] , 
        \R_DATA_TEMPR2[15] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR4[15] , 
        \R_DATA_TEMPR5[15] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR7[15] , 
        \R_DATA_TEMPR8[15] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR10[15] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR12[15] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR14[15] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR16[15] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR18[15] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR20[15] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR22[15] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR24[15] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR26[15] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR28[15] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR30[15] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR0[16] , \R_DATA_TEMPR1[16] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR3[16] , \R_DATA_TEMPR4[16] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR6[16] , \R_DATA_TEMPR7[16] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR9[16] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR11[16] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR13[16] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR15[16] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR17[16] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR19[16] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR21[16] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR23[16] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR25[16] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR27[16] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR29[16] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR31[16] , \R_DATA_TEMPR0[17] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR2[17] , \R_DATA_TEMPR3[17] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR5[17] , \R_DATA_TEMPR6[17] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR8[17] , \R_DATA_TEMPR9[17] , \R_DATA_TEMPR10[17] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR12[17] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR14[17] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR16[17] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR18[17] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR20[17] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR22[17] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR24[17] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR26[17] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR28[17] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR30[17] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR1[18] , 
        \R_DATA_TEMPR2[18] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR4[18] , 
        \R_DATA_TEMPR5[18] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR7[18] , 
        \R_DATA_TEMPR8[18] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR11[18] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR13[18] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR15[18] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR17[18] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR19[18] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR21[18] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR23[18] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR25[18] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR27[18] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR29[18] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR31[18] , \R_DATA_TEMPR0[19] , \R_DATA_TEMPR1[19] , 
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR3[19] , \R_DATA_TEMPR4[19] , 
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR6[19] , \R_DATA_TEMPR7[19] , 
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR9[19] , \R_DATA_TEMPR10[19] , 
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR12[19] , 
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR14[19] , 
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR16[19] , 
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR18[19] , 
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR20[19] , 
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR22[19] , 
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR24[19] , 
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR26[19] , 
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR28[19] , 
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR30[19] , 
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR0[20] , \R_DATA_TEMPR1[20] , 
        \R_DATA_TEMPR2[20] , \R_DATA_TEMPR3[20] , \R_DATA_TEMPR4[20] , 
        \R_DATA_TEMPR5[20] , \R_DATA_TEMPR6[20] , \R_DATA_TEMPR7[20] , 
        \R_DATA_TEMPR8[20] , \R_DATA_TEMPR9[20] , \R_DATA_TEMPR10[20] , 
        \R_DATA_TEMPR11[20] , \R_DATA_TEMPR12[20] , 
        \R_DATA_TEMPR13[20] , \R_DATA_TEMPR14[20] , 
        \R_DATA_TEMPR15[20] , \R_DATA_TEMPR16[20] , 
        \R_DATA_TEMPR17[20] , \R_DATA_TEMPR18[20] , 
        \R_DATA_TEMPR19[20] , \R_DATA_TEMPR20[20] , 
        \R_DATA_TEMPR21[20] , \R_DATA_TEMPR22[20] , 
        \R_DATA_TEMPR23[20] , \R_DATA_TEMPR24[20] , 
        \R_DATA_TEMPR25[20] , \R_DATA_TEMPR26[20] , 
        \R_DATA_TEMPR27[20] , \R_DATA_TEMPR28[20] , 
        \R_DATA_TEMPR29[20] , \R_DATA_TEMPR30[20] , 
        \R_DATA_TEMPR31[20] , \R_DATA_TEMPR0[21] , \R_DATA_TEMPR1[21] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR3[21] , \R_DATA_TEMPR4[21] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR6[21] , \R_DATA_TEMPR7[21] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR9[21] , \R_DATA_TEMPR10[21] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR12[21] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR14[21] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR16[21] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR18[21] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR20[21] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR22[21] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR24[21] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR26[21] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR28[21] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR30[21] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR0[22] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR2[22] , \R_DATA_TEMPR3[22] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR5[22] , \R_DATA_TEMPR6[22] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR8[22] , \R_DATA_TEMPR9[22] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR11[22] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR13[22] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR15[22] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR17[22] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR19[22] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR21[22] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR23[22] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR25[22] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR27[22] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR29[22] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR31[22] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR1[23] , 
        \R_DATA_TEMPR2[23] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR4[23] , 
        \R_DATA_TEMPR5[23] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR7[23] , 
        \R_DATA_TEMPR8[23] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR10[23] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR12[23] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR14[23] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR16[23] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR18[23] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR20[23] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR22[23] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR24[23] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR26[23] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR28[23] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR30[23] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR0[24] , \R_DATA_TEMPR1[24] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR3[24] , \R_DATA_TEMPR4[24] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR6[24] , \R_DATA_TEMPR7[24] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR9[24] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR11[24] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR13[24] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR15[24] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR17[24] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR19[24] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR21[24] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR23[24] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR25[24] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR27[24] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR29[24] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR31[24] , \R_DATA_TEMPR0[25] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR2[25] , \R_DATA_TEMPR3[25] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR5[25] , \R_DATA_TEMPR6[25] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR8[25] , \R_DATA_TEMPR9[25] , \R_DATA_TEMPR10[25] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR12[25] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR14[25] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR16[25] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR18[25] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR20[25] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR22[25] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR24[25] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR26[25] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR28[25] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR30[25] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR1[26] , 
        \R_DATA_TEMPR2[26] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR4[26] , 
        \R_DATA_TEMPR5[26] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR7[26] , 
        \R_DATA_TEMPR8[26] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR11[26] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR13[26] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR15[26] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR17[26] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR19[26] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR21[26] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR23[26] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR25[26] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR27[26] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR29[26] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR31[26] , \R_DATA_TEMPR0[27] , \R_DATA_TEMPR1[27] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR3[27] , \R_DATA_TEMPR4[27] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR6[27] , \R_DATA_TEMPR7[27] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR9[27] , \R_DATA_TEMPR10[27] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR12[27] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR14[27] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR16[27] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR18[27] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR20[27] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR22[27] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR24[27] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR26[27] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR28[27] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR30[27] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR0[28] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR2[28] , \R_DATA_TEMPR3[28] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR5[28] , \R_DATA_TEMPR6[28] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR8[28] , \R_DATA_TEMPR9[28] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR11[28] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR13[28] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR15[28] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR17[28] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR19[28] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR21[28] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR23[28] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR25[28] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR27[28] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR29[28] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR31[28] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR1[29] , 
        \R_DATA_TEMPR2[29] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR4[29] , 
        \R_DATA_TEMPR5[29] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR7[29] , 
        \R_DATA_TEMPR8[29] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR10[29] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR12[29] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR14[29] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR16[29] , 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR18[29] , 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR20[29] , 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR22[29] , 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR24[29] , 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR26[29] , 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR28[29] , 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR30[29] , 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR0[30] , \R_DATA_TEMPR1[30] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR3[30] , \R_DATA_TEMPR4[30] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR6[30] , \R_DATA_TEMPR7[30] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR9[30] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR11[30] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR13[30] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR15[30] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR17[30] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR19[30] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR21[30] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR23[30] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR25[30] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR27[30] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR29[30] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR31[30] , \R_DATA_TEMPR0[31] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR2[31] , \R_DATA_TEMPR3[31] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR5[31] , \R_DATA_TEMPR6[31] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR8[31] , \R_DATA_TEMPR9[31] , \R_DATA_TEMPR10[31] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR12[31] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR14[31] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR16[31] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR18[31] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR20[31] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR22[31] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR24[31] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR26[31] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR28[31] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR30[31] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR1[32] , 
        \R_DATA_TEMPR2[32] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR4[32] , 
        \R_DATA_TEMPR5[32] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR7[32] , 
        \R_DATA_TEMPR8[32] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR11[32] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR13[32] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR15[32] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR17[32] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR19[32] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR21[32] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR23[32] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR25[32] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR27[32] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR29[32] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR31[32] , \R_DATA_TEMPR0[33] , \R_DATA_TEMPR1[33] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR3[33] , \R_DATA_TEMPR4[33] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR6[33] , \R_DATA_TEMPR7[33] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR9[33] , \R_DATA_TEMPR10[33] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR12[33] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR14[33] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR16[33] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR18[33] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR20[33] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR22[33] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR24[33] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR26[33] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR28[33] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR30[33] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR0[34] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR2[34] , \R_DATA_TEMPR3[34] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR5[34] , \R_DATA_TEMPR6[34] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR8[34] , \R_DATA_TEMPR9[34] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR11[34] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR13[34] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR15[34] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR17[34] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR19[34] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR21[34] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR23[34] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR25[34] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR27[34] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR29[34] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR31[34] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR1[35] , 
        \R_DATA_TEMPR2[35] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR4[35] , 
        \R_DATA_TEMPR5[35] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR7[35] , 
        \R_DATA_TEMPR8[35] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR10[35] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR12[35] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR14[35] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR16[35] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR18[35] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR20[35] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR22[35] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR24[35] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR26[35] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR28[35] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR30[35] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR0[36] , \R_DATA_TEMPR1[36] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR3[36] , \R_DATA_TEMPR4[36] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR6[36] , \R_DATA_TEMPR7[36] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR9[36] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR11[36] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR13[36] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR15[36] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR17[36] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR19[36] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR21[36] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR23[36] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR25[36] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR27[36] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR29[36] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR31[36] , \R_DATA_TEMPR0[37] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR2[37] , \R_DATA_TEMPR3[37] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR5[37] , \R_DATA_TEMPR6[37] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR8[37] , \R_DATA_TEMPR9[37] , \R_DATA_TEMPR10[37] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR12[37] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR14[37] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR16[37] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR18[37] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR20[37] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR22[37] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR24[37] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR26[37] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR28[37] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR30[37] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR1[38] , 
        \R_DATA_TEMPR2[38] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR4[38] , 
        \R_DATA_TEMPR5[38] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR7[38] , 
        \R_DATA_TEMPR8[38] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR11[38] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR13[38] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR15[38] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR17[38] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR19[38] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR21[38] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR23[38] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR25[38] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR27[38] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR29[38] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR31[38] , \R_DATA_TEMPR0[39] , \R_DATA_TEMPR1[39] , 
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR3[39] , \R_DATA_TEMPR4[39] , 
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR6[39] , \R_DATA_TEMPR7[39] , 
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR9[39] , \R_DATA_TEMPR10[39] , 
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR12[39] , 
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR14[39] , 
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR16[39] , 
        \R_DATA_TEMPR17[39] , \R_DATA_TEMPR18[39] , 
        \R_DATA_TEMPR19[39] , \R_DATA_TEMPR20[39] , 
        \R_DATA_TEMPR21[39] , \R_DATA_TEMPR22[39] , 
        \R_DATA_TEMPR23[39] , \R_DATA_TEMPR24[39] , 
        \R_DATA_TEMPR25[39] , \R_DATA_TEMPR26[39] , 
        \R_DATA_TEMPR27[39] , \R_DATA_TEMPR28[39] , 
        \R_DATA_TEMPR29[39] , \R_DATA_TEMPR30[39] , 
        \R_DATA_TEMPR31[39] , \BLKX0[0] , \BLKY0[0] , \BLKX1[0] , 
        \BLKY1[0] , \BLKX2[0] , \BLKX2[1] , \BLKX2[2] , \BLKX2[3] , 
        \BLKX2[4] , \BLKX2[5] , \BLKX2[6] , \BLKX2[7] , \BLKY2[0] , 
        \BLKY2[1] , \BLKY2[2] , \BLKY2[3] , \BLKY2[4] , \BLKY2[5] , 
        \BLKY2[6] , \BLKY2[7] , \ACCESS_BUSY[0][0] , 
        \SB_CORRECT[0][0] , \DB_DETECT[0][0] , \ACCESS_BUSY[0][1] , 
        \SB_CORRECT[0][1] , \DB_DETECT[0][1] , \ACCESS_BUSY[0][2] , 
        \SB_CORRECT[0][2] , \DB_DETECT[0][2] , \ACCESS_BUSY[0][3] , 
        \SB_CORRECT[0][3] , \DB_DETECT[0][3] , \ACCESS_BUSY[0][4] , 
        \SB_CORRECT[0][4] , \DB_DETECT[0][4] , \ACCESS_BUSY[0][5] , 
        \SB_CORRECT[0][5] , \DB_DETECT[0][5] , \ACCESS_BUSY[0][6] , 
        \SB_CORRECT[0][6] , \DB_DETECT[0][6] , \ACCESS_BUSY[0][7] , 
        \SB_CORRECT[0][7] , \DB_DETECT[0][7] , \ACCESS_BUSY[0][8] , 
        \SB_CORRECT[0][8] , \DB_DETECT[0][8] , \ACCESS_BUSY[0][9] , 
        \SB_CORRECT[0][9] , \DB_DETECT[0][9] , \ACCESS_BUSY[0][10] , 
        \SB_CORRECT[0][10] , \DB_DETECT[0][10] , \ACCESS_BUSY[0][11] , 
        \SB_CORRECT[0][11] , \DB_DETECT[0][11] , \ACCESS_BUSY[0][12] , 
        \SB_CORRECT[0][12] , \DB_DETECT[0][12] , \ACCESS_BUSY[0][13] , 
        \SB_CORRECT[0][13] , \DB_DETECT[0][13] , \ACCESS_BUSY[0][14] , 
        \SB_CORRECT[0][14] , \DB_DETECT[0][14] , \ACCESS_BUSY[0][15] , 
        \SB_CORRECT[0][15] , \DB_DETECT[0][15] , \ACCESS_BUSY[0][16] , 
        \SB_CORRECT[0][16] , \DB_DETECT[0][16] , \ACCESS_BUSY[0][17] , 
        \SB_CORRECT[0][17] , \DB_DETECT[0][17] , \ACCESS_BUSY[0][18] , 
        \SB_CORRECT[0][18] , \DB_DETECT[0][18] , \ACCESS_BUSY[0][19] , 
        \SB_CORRECT[0][19] , \DB_DETECT[0][19] , \ACCESS_BUSY[1][0] , 
        \SB_CORRECT[1][0] , \DB_DETECT[1][0] , \ACCESS_BUSY[1][1] , 
        \SB_CORRECT[1][1] , \DB_DETECT[1][1] , \ACCESS_BUSY[1][2] , 
        \SB_CORRECT[1][2] , \DB_DETECT[1][2] , \ACCESS_BUSY[1][3] , 
        \SB_CORRECT[1][3] , \DB_DETECT[1][3] , \ACCESS_BUSY[1][4] , 
        \SB_CORRECT[1][4] , \DB_DETECT[1][4] , \ACCESS_BUSY[1][5] , 
        \SB_CORRECT[1][5] , \DB_DETECT[1][5] , \ACCESS_BUSY[1][6] , 
        \SB_CORRECT[1][6] , \DB_DETECT[1][6] , \ACCESS_BUSY[1][7] , 
        \SB_CORRECT[1][7] , \DB_DETECT[1][7] , \ACCESS_BUSY[1][8] , 
        \SB_CORRECT[1][8] , \DB_DETECT[1][8] , \ACCESS_BUSY[1][9] , 
        \SB_CORRECT[1][9] , \DB_DETECT[1][9] , \ACCESS_BUSY[1][10] , 
        \SB_CORRECT[1][10] , \DB_DETECT[1][10] , \ACCESS_BUSY[1][11] , 
        \SB_CORRECT[1][11] , \DB_DETECT[1][11] , \ACCESS_BUSY[1][12] , 
        \SB_CORRECT[1][12] , \DB_DETECT[1][12] , \ACCESS_BUSY[1][13] , 
        \SB_CORRECT[1][13] , \DB_DETECT[1][13] , \ACCESS_BUSY[1][14] , 
        \SB_CORRECT[1][14] , \DB_DETECT[1][14] , \ACCESS_BUSY[1][15] , 
        \SB_CORRECT[1][15] , \DB_DETECT[1][15] , \ACCESS_BUSY[1][16] , 
        \SB_CORRECT[1][16] , \DB_DETECT[1][16] , \ACCESS_BUSY[1][17] , 
        \SB_CORRECT[1][17] , \DB_DETECT[1][17] , \ACCESS_BUSY[1][18] , 
        \SB_CORRECT[1][18] , \DB_DETECT[1][18] , \ACCESS_BUSY[1][19] , 
        \SB_CORRECT[1][19] , \DB_DETECT[1][19] , \ACCESS_BUSY[2][0] , 
        \SB_CORRECT[2][0] , \DB_DETECT[2][0] , \ACCESS_BUSY[2][1] , 
        \SB_CORRECT[2][1] , \DB_DETECT[2][1] , \ACCESS_BUSY[2][2] , 
        \SB_CORRECT[2][2] , \DB_DETECT[2][2] , \ACCESS_BUSY[2][3] , 
        \SB_CORRECT[2][3] , \DB_DETECT[2][3] , \ACCESS_BUSY[2][4] , 
        \SB_CORRECT[2][4] , \DB_DETECT[2][4] , \ACCESS_BUSY[2][5] , 
        \SB_CORRECT[2][5] , \DB_DETECT[2][5] , \ACCESS_BUSY[2][6] , 
        \SB_CORRECT[2][6] , \DB_DETECT[2][6] , \ACCESS_BUSY[2][7] , 
        \SB_CORRECT[2][7] , \DB_DETECT[2][7] , \ACCESS_BUSY[2][8] , 
        \SB_CORRECT[2][8] , \DB_DETECT[2][8] , \ACCESS_BUSY[2][9] , 
        \SB_CORRECT[2][9] , \DB_DETECT[2][9] , \ACCESS_BUSY[2][10] , 
        \SB_CORRECT[2][10] , \DB_DETECT[2][10] , \ACCESS_BUSY[2][11] , 
        \SB_CORRECT[2][11] , \DB_DETECT[2][11] , \ACCESS_BUSY[2][12] , 
        \SB_CORRECT[2][12] , \DB_DETECT[2][12] , \ACCESS_BUSY[2][13] , 
        \SB_CORRECT[2][13] , \DB_DETECT[2][13] , \ACCESS_BUSY[2][14] , 
        \SB_CORRECT[2][14] , \DB_DETECT[2][14] , \ACCESS_BUSY[2][15] , 
        \SB_CORRECT[2][15] , \DB_DETECT[2][15] , \ACCESS_BUSY[2][16] , 
        \SB_CORRECT[2][16] , \DB_DETECT[2][16] , \ACCESS_BUSY[2][17] , 
        \SB_CORRECT[2][17] , \DB_DETECT[2][17] , \ACCESS_BUSY[2][18] , 
        \SB_CORRECT[2][18] , \DB_DETECT[2][18] , \ACCESS_BUSY[2][19] , 
        \SB_CORRECT[2][19] , \DB_DETECT[2][19] , \ACCESS_BUSY[3][0] , 
        \SB_CORRECT[3][0] , \DB_DETECT[3][0] , \ACCESS_BUSY[3][1] , 
        \SB_CORRECT[3][1] , \DB_DETECT[3][1] , \ACCESS_BUSY[3][2] , 
        \SB_CORRECT[3][2] , \DB_DETECT[3][2] , \ACCESS_BUSY[3][3] , 
        \SB_CORRECT[3][3] , \DB_DETECT[3][3] , \ACCESS_BUSY[3][4] , 
        \SB_CORRECT[3][4] , \DB_DETECT[3][4] , \ACCESS_BUSY[3][5] , 
        \SB_CORRECT[3][5] , \DB_DETECT[3][5] , \ACCESS_BUSY[3][6] , 
        \SB_CORRECT[3][6] , \DB_DETECT[3][6] , \ACCESS_BUSY[3][7] , 
        \SB_CORRECT[3][7] , \DB_DETECT[3][7] , \ACCESS_BUSY[3][8] , 
        \SB_CORRECT[3][8] , \DB_DETECT[3][8] , \ACCESS_BUSY[3][9] , 
        \SB_CORRECT[3][9] , \DB_DETECT[3][9] , \ACCESS_BUSY[3][10] , 
        \SB_CORRECT[3][10] , \DB_DETECT[3][10] , \ACCESS_BUSY[3][11] , 
        \SB_CORRECT[3][11] , \DB_DETECT[3][11] , \ACCESS_BUSY[3][12] , 
        \SB_CORRECT[3][12] , \DB_DETECT[3][12] , \ACCESS_BUSY[3][13] , 
        \SB_CORRECT[3][13] , \DB_DETECT[3][13] , \ACCESS_BUSY[3][14] , 
        \SB_CORRECT[3][14] , \DB_DETECT[3][14] , \ACCESS_BUSY[3][15] , 
        \SB_CORRECT[3][15] , \DB_DETECT[3][15] , \ACCESS_BUSY[3][16] , 
        \SB_CORRECT[3][16] , \DB_DETECT[3][16] , \ACCESS_BUSY[3][17] , 
        \SB_CORRECT[3][17] , \DB_DETECT[3][17] , \ACCESS_BUSY[3][18] , 
        \SB_CORRECT[3][18] , \DB_DETECT[3][18] , \ACCESS_BUSY[3][19] , 
        \SB_CORRECT[3][19] , \DB_DETECT[3][19] , \ACCESS_BUSY[4][0] , 
        \SB_CORRECT[4][0] , \DB_DETECT[4][0] , \ACCESS_BUSY[4][1] , 
        \SB_CORRECT[4][1] , \DB_DETECT[4][1] , \ACCESS_BUSY[4][2] , 
        \SB_CORRECT[4][2] , \DB_DETECT[4][2] , \ACCESS_BUSY[4][3] , 
        \SB_CORRECT[4][3] , \DB_DETECT[4][3] , \ACCESS_BUSY[4][4] , 
        \SB_CORRECT[4][4] , \DB_DETECT[4][4] , \ACCESS_BUSY[4][5] , 
        \SB_CORRECT[4][5] , \DB_DETECT[4][5] , \ACCESS_BUSY[4][6] , 
        \SB_CORRECT[4][6] , \DB_DETECT[4][6] , \ACCESS_BUSY[4][7] , 
        \SB_CORRECT[4][7] , \DB_DETECT[4][7] , \ACCESS_BUSY[4][8] , 
        \SB_CORRECT[4][8] , \DB_DETECT[4][8] , \ACCESS_BUSY[4][9] , 
        \SB_CORRECT[4][9] , \DB_DETECT[4][9] , \ACCESS_BUSY[4][10] , 
        \SB_CORRECT[4][10] , \DB_DETECT[4][10] , \ACCESS_BUSY[4][11] , 
        \SB_CORRECT[4][11] , \DB_DETECT[4][11] , \ACCESS_BUSY[4][12] , 
        \SB_CORRECT[4][12] , \DB_DETECT[4][12] , \ACCESS_BUSY[4][13] , 
        \SB_CORRECT[4][13] , \DB_DETECT[4][13] , \ACCESS_BUSY[4][14] , 
        \SB_CORRECT[4][14] , \DB_DETECT[4][14] , \ACCESS_BUSY[4][15] , 
        \SB_CORRECT[4][15] , \DB_DETECT[4][15] , \ACCESS_BUSY[4][16] , 
        \SB_CORRECT[4][16] , \DB_DETECT[4][16] , \ACCESS_BUSY[4][17] , 
        \SB_CORRECT[4][17] , \DB_DETECT[4][17] , \ACCESS_BUSY[4][18] , 
        \SB_CORRECT[4][18] , \DB_DETECT[4][18] , \ACCESS_BUSY[4][19] , 
        \SB_CORRECT[4][19] , \DB_DETECT[4][19] , \ACCESS_BUSY[5][0] , 
        \SB_CORRECT[5][0] , \DB_DETECT[5][0] , \ACCESS_BUSY[5][1] , 
        \SB_CORRECT[5][1] , \DB_DETECT[5][1] , \ACCESS_BUSY[5][2] , 
        \SB_CORRECT[5][2] , \DB_DETECT[5][2] , \ACCESS_BUSY[5][3] , 
        \SB_CORRECT[5][3] , \DB_DETECT[5][3] , \ACCESS_BUSY[5][4] , 
        \SB_CORRECT[5][4] , \DB_DETECT[5][4] , \ACCESS_BUSY[5][5] , 
        \SB_CORRECT[5][5] , \DB_DETECT[5][5] , \ACCESS_BUSY[5][6] , 
        \SB_CORRECT[5][6] , \DB_DETECT[5][6] , \ACCESS_BUSY[5][7] , 
        \SB_CORRECT[5][7] , \DB_DETECT[5][7] , \ACCESS_BUSY[5][8] , 
        \SB_CORRECT[5][8] , \DB_DETECT[5][8] , \ACCESS_BUSY[5][9] , 
        \SB_CORRECT[5][9] , \DB_DETECT[5][9] , \ACCESS_BUSY[5][10] , 
        \SB_CORRECT[5][10] , \DB_DETECT[5][10] , \ACCESS_BUSY[5][11] , 
        \SB_CORRECT[5][11] , \DB_DETECT[5][11] , \ACCESS_BUSY[5][12] , 
        \SB_CORRECT[5][12] , \DB_DETECT[5][12] , \ACCESS_BUSY[5][13] , 
        \SB_CORRECT[5][13] , \DB_DETECT[5][13] , \ACCESS_BUSY[5][14] , 
        \SB_CORRECT[5][14] , \DB_DETECT[5][14] , \ACCESS_BUSY[5][15] , 
        \SB_CORRECT[5][15] , \DB_DETECT[5][15] , \ACCESS_BUSY[5][16] , 
        \SB_CORRECT[5][16] , \DB_DETECT[5][16] , \ACCESS_BUSY[5][17] , 
        \SB_CORRECT[5][17] , \DB_DETECT[5][17] , \ACCESS_BUSY[5][18] , 
        \SB_CORRECT[5][18] , \DB_DETECT[5][18] , \ACCESS_BUSY[5][19] , 
        \SB_CORRECT[5][19] , \DB_DETECT[5][19] , \ACCESS_BUSY[6][0] , 
        \SB_CORRECT[6][0] , \DB_DETECT[6][0] , \ACCESS_BUSY[6][1] , 
        \SB_CORRECT[6][1] , \DB_DETECT[6][1] , \ACCESS_BUSY[6][2] , 
        \SB_CORRECT[6][2] , \DB_DETECT[6][2] , \ACCESS_BUSY[6][3] , 
        \SB_CORRECT[6][3] , \DB_DETECT[6][3] , \ACCESS_BUSY[6][4] , 
        \SB_CORRECT[6][4] , \DB_DETECT[6][4] , \ACCESS_BUSY[6][5] , 
        \SB_CORRECT[6][5] , \DB_DETECT[6][5] , \ACCESS_BUSY[6][6] , 
        \SB_CORRECT[6][6] , \DB_DETECT[6][6] , \ACCESS_BUSY[6][7] , 
        \SB_CORRECT[6][7] , \DB_DETECT[6][7] , \ACCESS_BUSY[6][8] , 
        \SB_CORRECT[6][8] , \DB_DETECT[6][8] , \ACCESS_BUSY[6][9] , 
        \SB_CORRECT[6][9] , \DB_DETECT[6][9] , \ACCESS_BUSY[6][10] , 
        \SB_CORRECT[6][10] , \DB_DETECT[6][10] , \ACCESS_BUSY[6][11] , 
        \SB_CORRECT[6][11] , \DB_DETECT[6][11] , \ACCESS_BUSY[6][12] , 
        \SB_CORRECT[6][12] , \DB_DETECT[6][12] , \ACCESS_BUSY[6][13] , 
        \SB_CORRECT[6][13] , \DB_DETECT[6][13] , \ACCESS_BUSY[6][14] , 
        \SB_CORRECT[6][14] , \DB_DETECT[6][14] , \ACCESS_BUSY[6][15] , 
        \SB_CORRECT[6][15] , \DB_DETECT[6][15] , \ACCESS_BUSY[6][16] , 
        \SB_CORRECT[6][16] , \DB_DETECT[6][16] , \ACCESS_BUSY[6][17] , 
        \SB_CORRECT[6][17] , \DB_DETECT[6][17] , \ACCESS_BUSY[6][18] , 
        \SB_CORRECT[6][18] , \DB_DETECT[6][18] , \ACCESS_BUSY[6][19] , 
        \SB_CORRECT[6][19] , \DB_DETECT[6][19] , \ACCESS_BUSY[7][0] , 
        \SB_CORRECT[7][0] , \DB_DETECT[7][0] , \ACCESS_BUSY[7][1] , 
        \SB_CORRECT[7][1] , \DB_DETECT[7][1] , \ACCESS_BUSY[7][2] , 
        \SB_CORRECT[7][2] , \DB_DETECT[7][2] , \ACCESS_BUSY[7][3] , 
        \SB_CORRECT[7][3] , \DB_DETECT[7][3] , \ACCESS_BUSY[7][4] , 
        \SB_CORRECT[7][4] , \DB_DETECT[7][4] , \ACCESS_BUSY[7][5] , 
        \SB_CORRECT[7][5] , \DB_DETECT[7][5] , \ACCESS_BUSY[7][6] , 
        \SB_CORRECT[7][6] , \DB_DETECT[7][6] , \ACCESS_BUSY[7][7] , 
        \SB_CORRECT[7][7] , \DB_DETECT[7][7] , \ACCESS_BUSY[7][8] , 
        \SB_CORRECT[7][8] , \DB_DETECT[7][8] , \ACCESS_BUSY[7][9] , 
        \SB_CORRECT[7][9] , \DB_DETECT[7][9] , \ACCESS_BUSY[7][10] , 
        \SB_CORRECT[7][10] , \DB_DETECT[7][10] , \ACCESS_BUSY[7][11] , 
        \SB_CORRECT[7][11] , \DB_DETECT[7][11] , \ACCESS_BUSY[7][12] , 
        \SB_CORRECT[7][12] , \DB_DETECT[7][12] , \ACCESS_BUSY[7][13] , 
        \SB_CORRECT[7][13] , \DB_DETECT[7][13] , \ACCESS_BUSY[7][14] , 
        \SB_CORRECT[7][14] , \DB_DETECT[7][14] , \ACCESS_BUSY[7][15] , 
        \SB_CORRECT[7][15] , \DB_DETECT[7][15] , \ACCESS_BUSY[7][16] , 
        \SB_CORRECT[7][16] , \DB_DETECT[7][16] , \ACCESS_BUSY[7][17] , 
        \SB_CORRECT[7][17] , \DB_DETECT[7][17] , \ACCESS_BUSY[7][18] , 
        \SB_CORRECT[7][18] , \DB_DETECT[7][18] , \ACCESS_BUSY[7][19] , 
        \SB_CORRECT[7][19] , \DB_DETECT[7][19] , \ACCESS_BUSY[8][0] , 
        \SB_CORRECT[8][0] , \DB_DETECT[8][0] , \ACCESS_BUSY[8][1] , 
        \SB_CORRECT[8][1] , \DB_DETECT[8][1] , \ACCESS_BUSY[8][2] , 
        \SB_CORRECT[8][2] , \DB_DETECT[8][2] , \ACCESS_BUSY[8][3] , 
        \SB_CORRECT[8][3] , \DB_DETECT[8][3] , \ACCESS_BUSY[8][4] , 
        \SB_CORRECT[8][4] , \DB_DETECT[8][4] , \ACCESS_BUSY[8][5] , 
        \SB_CORRECT[8][5] , \DB_DETECT[8][5] , \ACCESS_BUSY[8][6] , 
        \SB_CORRECT[8][6] , \DB_DETECT[8][6] , \ACCESS_BUSY[8][7] , 
        \SB_CORRECT[8][7] , \DB_DETECT[8][7] , \ACCESS_BUSY[8][8] , 
        \SB_CORRECT[8][8] , \DB_DETECT[8][8] , \ACCESS_BUSY[8][9] , 
        \SB_CORRECT[8][9] , \DB_DETECT[8][9] , \ACCESS_BUSY[8][10] , 
        \SB_CORRECT[8][10] , \DB_DETECT[8][10] , \ACCESS_BUSY[8][11] , 
        \SB_CORRECT[8][11] , \DB_DETECT[8][11] , \ACCESS_BUSY[8][12] , 
        \SB_CORRECT[8][12] , \DB_DETECT[8][12] , \ACCESS_BUSY[8][13] , 
        \SB_CORRECT[8][13] , \DB_DETECT[8][13] , \ACCESS_BUSY[8][14] , 
        \SB_CORRECT[8][14] , \DB_DETECT[8][14] , \ACCESS_BUSY[8][15] , 
        \SB_CORRECT[8][15] , \DB_DETECT[8][15] , \ACCESS_BUSY[8][16] , 
        \SB_CORRECT[8][16] , \DB_DETECT[8][16] , \ACCESS_BUSY[8][17] , 
        \SB_CORRECT[8][17] , \DB_DETECT[8][17] , \ACCESS_BUSY[8][18] , 
        \SB_CORRECT[8][18] , \DB_DETECT[8][18] , \ACCESS_BUSY[8][19] , 
        \SB_CORRECT[8][19] , \DB_DETECT[8][19] , \ACCESS_BUSY[9][0] , 
        \SB_CORRECT[9][0] , \DB_DETECT[9][0] , \ACCESS_BUSY[9][1] , 
        \SB_CORRECT[9][1] , \DB_DETECT[9][1] , \ACCESS_BUSY[9][2] , 
        \SB_CORRECT[9][2] , \DB_DETECT[9][2] , \ACCESS_BUSY[9][3] , 
        \SB_CORRECT[9][3] , \DB_DETECT[9][3] , \ACCESS_BUSY[9][4] , 
        \SB_CORRECT[9][4] , \DB_DETECT[9][4] , \ACCESS_BUSY[9][5] , 
        \SB_CORRECT[9][5] , \DB_DETECT[9][5] , \ACCESS_BUSY[9][6] , 
        \SB_CORRECT[9][6] , \DB_DETECT[9][6] , \ACCESS_BUSY[9][7] , 
        \SB_CORRECT[9][7] , \DB_DETECT[9][7] , \ACCESS_BUSY[9][8] , 
        \SB_CORRECT[9][8] , \DB_DETECT[9][8] , \ACCESS_BUSY[9][9] , 
        \SB_CORRECT[9][9] , \DB_DETECT[9][9] , \ACCESS_BUSY[9][10] , 
        \SB_CORRECT[9][10] , \DB_DETECT[9][10] , \ACCESS_BUSY[9][11] , 
        \SB_CORRECT[9][11] , \DB_DETECT[9][11] , \ACCESS_BUSY[9][12] , 
        \SB_CORRECT[9][12] , \DB_DETECT[9][12] , \ACCESS_BUSY[9][13] , 
        \SB_CORRECT[9][13] , \DB_DETECT[9][13] , \ACCESS_BUSY[9][14] , 
        \SB_CORRECT[9][14] , \DB_DETECT[9][14] , \ACCESS_BUSY[9][15] , 
        \SB_CORRECT[9][15] , \DB_DETECT[9][15] , \ACCESS_BUSY[9][16] , 
        \SB_CORRECT[9][16] , \DB_DETECT[9][16] , \ACCESS_BUSY[9][17] , 
        \SB_CORRECT[9][17] , \DB_DETECT[9][17] , \ACCESS_BUSY[9][18] , 
        \SB_CORRECT[9][18] , \DB_DETECT[9][18] , \ACCESS_BUSY[9][19] , 
        \SB_CORRECT[9][19] , \DB_DETECT[9][19] , \ACCESS_BUSY[10][0] , 
        \SB_CORRECT[10][0] , \DB_DETECT[10][0] , \ACCESS_BUSY[10][1] , 
        \SB_CORRECT[10][1] , \DB_DETECT[10][1] , \ACCESS_BUSY[10][2] , 
        \SB_CORRECT[10][2] , \DB_DETECT[10][2] , \ACCESS_BUSY[10][3] , 
        \SB_CORRECT[10][3] , \DB_DETECT[10][3] , \ACCESS_BUSY[10][4] , 
        \SB_CORRECT[10][4] , \DB_DETECT[10][4] , \ACCESS_BUSY[10][5] , 
        \SB_CORRECT[10][5] , \DB_DETECT[10][5] , \ACCESS_BUSY[10][6] , 
        \SB_CORRECT[10][6] , \DB_DETECT[10][6] , \ACCESS_BUSY[10][7] , 
        \SB_CORRECT[10][7] , \DB_DETECT[10][7] , \ACCESS_BUSY[10][8] , 
        \SB_CORRECT[10][8] , \DB_DETECT[10][8] , \ACCESS_BUSY[10][9] , 
        \SB_CORRECT[10][9] , \DB_DETECT[10][9] , \ACCESS_BUSY[10][10] , 
        \SB_CORRECT[10][10] , \DB_DETECT[10][10] , 
        \ACCESS_BUSY[10][11] , \SB_CORRECT[10][11] , 
        \DB_DETECT[10][11] , \ACCESS_BUSY[10][12] , 
        \SB_CORRECT[10][12] , \DB_DETECT[10][12] , 
        \ACCESS_BUSY[10][13] , \SB_CORRECT[10][13] , 
        \DB_DETECT[10][13] , \ACCESS_BUSY[10][14] , 
        \SB_CORRECT[10][14] , \DB_DETECT[10][14] , 
        \ACCESS_BUSY[10][15] , \SB_CORRECT[10][15] , 
        \DB_DETECT[10][15] , \ACCESS_BUSY[10][16] , 
        \SB_CORRECT[10][16] , \DB_DETECT[10][16] , 
        \ACCESS_BUSY[10][17] , \SB_CORRECT[10][17] , 
        \DB_DETECT[10][17] , \ACCESS_BUSY[10][18] , 
        \SB_CORRECT[10][18] , \DB_DETECT[10][18] , 
        \ACCESS_BUSY[10][19] , \SB_CORRECT[10][19] , 
        \DB_DETECT[10][19] , \ACCESS_BUSY[11][0] , \SB_CORRECT[11][0] , 
        \DB_DETECT[11][0] , \ACCESS_BUSY[11][1] , \SB_CORRECT[11][1] , 
        \DB_DETECT[11][1] , \ACCESS_BUSY[11][2] , \SB_CORRECT[11][2] , 
        \DB_DETECT[11][2] , \ACCESS_BUSY[11][3] , \SB_CORRECT[11][3] , 
        \DB_DETECT[11][3] , \ACCESS_BUSY[11][4] , \SB_CORRECT[11][4] , 
        \DB_DETECT[11][4] , \ACCESS_BUSY[11][5] , \SB_CORRECT[11][5] , 
        \DB_DETECT[11][5] , \ACCESS_BUSY[11][6] , \SB_CORRECT[11][6] , 
        \DB_DETECT[11][6] , \ACCESS_BUSY[11][7] , \SB_CORRECT[11][7] , 
        \DB_DETECT[11][7] , \ACCESS_BUSY[11][8] , \SB_CORRECT[11][8] , 
        \DB_DETECT[11][8] , \ACCESS_BUSY[11][9] , \SB_CORRECT[11][9] , 
        \DB_DETECT[11][9] , \ACCESS_BUSY[11][10] , 
        \SB_CORRECT[11][10] , \DB_DETECT[11][10] , 
        \ACCESS_BUSY[11][11] , \SB_CORRECT[11][11] , 
        \DB_DETECT[11][11] , \ACCESS_BUSY[11][12] , 
        \SB_CORRECT[11][12] , \DB_DETECT[11][12] , 
        \ACCESS_BUSY[11][13] , \SB_CORRECT[11][13] , 
        \DB_DETECT[11][13] , \ACCESS_BUSY[11][14] , 
        \SB_CORRECT[11][14] , \DB_DETECT[11][14] , 
        \ACCESS_BUSY[11][15] , \SB_CORRECT[11][15] , 
        \DB_DETECT[11][15] , \ACCESS_BUSY[11][16] , 
        \SB_CORRECT[11][16] , \DB_DETECT[11][16] , 
        \ACCESS_BUSY[11][17] , \SB_CORRECT[11][17] , 
        \DB_DETECT[11][17] , \ACCESS_BUSY[11][18] , 
        \SB_CORRECT[11][18] , \DB_DETECT[11][18] , 
        \ACCESS_BUSY[11][19] , \SB_CORRECT[11][19] , 
        \DB_DETECT[11][19] , \ACCESS_BUSY[12][0] , \SB_CORRECT[12][0] , 
        \DB_DETECT[12][0] , \ACCESS_BUSY[12][1] , \SB_CORRECT[12][1] , 
        \DB_DETECT[12][1] , \ACCESS_BUSY[12][2] , \SB_CORRECT[12][2] , 
        \DB_DETECT[12][2] , \ACCESS_BUSY[12][3] , \SB_CORRECT[12][3] , 
        \DB_DETECT[12][3] , \ACCESS_BUSY[12][4] , \SB_CORRECT[12][4] , 
        \DB_DETECT[12][4] , \ACCESS_BUSY[12][5] , \SB_CORRECT[12][5] , 
        \DB_DETECT[12][5] , \ACCESS_BUSY[12][6] , \SB_CORRECT[12][6] , 
        \DB_DETECT[12][6] , \ACCESS_BUSY[12][7] , \SB_CORRECT[12][7] , 
        \DB_DETECT[12][7] , \ACCESS_BUSY[12][8] , \SB_CORRECT[12][8] , 
        \DB_DETECT[12][8] , \ACCESS_BUSY[12][9] , \SB_CORRECT[12][9] , 
        \DB_DETECT[12][9] , \ACCESS_BUSY[12][10] , 
        \SB_CORRECT[12][10] , \DB_DETECT[12][10] , 
        \ACCESS_BUSY[12][11] , \SB_CORRECT[12][11] , 
        \DB_DETECT[12][11] , \ACCESS_BUSY[12][12] , 
        \SB_CORRECT[12][12] , \DB_DETECT[12][12] , 
        \ACCESS_BUSY[12][13] , \SB_CORRECT[12][13] , 
        \DB_DETECT[12][13] , \ACCESS_BUSY[12][14] , 
        \SB_CORRECT[12][14] , \DB_DETECT[12][14] , 
        \ACCESS_BUSY[12][15] , \SB_CORRECT[12][15] , 
        \DB_DETECT[12][15] , \ACCESS_BUSY[12][16] , 
        \SB_CORRECT[12][16] , \DB_DETECT[12][16] , 
        \ACCESS_BUSY[12][17] , \SB_CORRECT[12][17] , 
        \DB_DETECT[12][17] , \ACCESS_BUSY[12][18] , 
        \SB_CORRECT[12][18] , \DB_DETECT[12][18] , 
        \ACCESS_BUSY[12][19] , \SB_CORRECT[12][19] , 
        \DB_DETECT[12][19] , \ACCESS_BUSY[13][0] , \SB_CORRECT[13][0] , 
        \DB_DETECT[13][0] , \ACCESS_BUSY[13][1] , \SB_CORRECT[13][1] , 
        \DB_DETECT[13][1] , \ACCESS_BUSY[13][2] , \SB_CORRECT[13][2] , 
        \DB_DETECT[13][2] , \ACCESS_BUSY[13][3] , \SB_CORRECT[13][3] , 
        \DB_DETECT[13][3] , \ACCESS_BUSY[13][4] , \SB_CORRECT[13][4] , 
        \DB_DETECT[13][4] , \ACCESS_BUSY[13][5] , \SB_CORRECT[13][5] , 
        \DB_DETECT[13][5] , \ACCESS_BUSY[13][6] , \SB_CORRECT[13][6] , 
        \DB_DETECT[13][6] , \ACCESS_BUSY[13][7] , \SB_CORRECT[13][7] , 
        \DB_DETECT[13][7] , \ACCESS_BUSY[13][8] , \SB_CORRECT[13][8] , 
        \DB_DETECT[13][8] , \ACCESS_BUSY[13][9] , \SB_CORRECT[13][9] , 
        \DB_DETECT[13][9] , \ACCESS_BUSY[13][10] , 
        \SB_CORRECT[13][10] , \DB_DETECT[13][10] , 
        \ACCESS_BUSY[13][11] , \SB_CORRECT[13][11] , 
        \DB_DETECT[13][11] , \ACCESS_BUSY[13][12] , 
        \SB_CORRECT[13][12] , \DB_DETECT[13][12] , 
        \ACCESS_BUSY[13][13] , \SB_CORRECT[13][13] , 
        \DB_DETECT[13][13] , \ACCESS_BUSY[13][14] , 
        \SB_CORRECT[13][14] , \DB_DETECT[13][14] , 
        \ACCESS_BUSY[13][15] , \SB_CORRECT[13][15] , 
        \DB_DETECT[13][15] , \ACCESS_BUSY[13][16] , 
        \SB_CORRECT[13][16] , \DB_DETECT[13][16] , 
        \ACCESS_BUSY[13][17] , \SB_CORRECT[13][17] , 
        \DB_DETECT[13][17] , \ACCESS_BUSY[13][18] , 
        \SB_CORRECT[13][18] , \DB_DETECT[13][18] , 
        \ACCESS_BUSY[13][19] , \SB_CORRECT[13][19] , 
        \DB_DETECT[13][19] , \ACCESS_BUSY[14][0] , \SB_CORRECT[14][0] , 
        \DB_DETECT[14][0] , \ACCESS_BUSY[14][1] , \SB_CORRECT[14][1] , 
        \DB_DETECT[14][1] , \ACCESS_BUSY[14][2] , \SB_CORRECT[14][2] , 
        \DB_DETECT[14][2] , \ACCESS_BUSY[14][3] , \SB_CORRECT[14][3] , 
        \DB_DETECT[14][3] , \ACCESS_BUSY[14][4] , \SB_CORRECT[14][4] , 
        \DB_DETECT[14][4] , \ACCESS_BUSY[14][5] , \SB_CORRECT[14][5] , 
        \DB_DETECT[14][5] , \ACCESS_BUSY[14][6] , \SB_CORRECT[14][6] , 
        \DB_DETECT[14][6] , \ACCESS_BUSY[14][7] , \SB_CORRECT[14][7] , 
        \DB_DETECT[14][7] , \ACCESS_BUSY[14][8] , \SB_CORRECT[14][8] , 
        \DB_DETECT[14][8] , \ACCESS_BUSY[14][9] , \SB_CORRECT[14][9] , 
        \DB_DETECT[14][9] , \ACCESS_BUSY[14][10] , 
        \SB_CORRECT[14][10] , \DB_DETECT[14][10] , 
        \ACCESS_BUSY[14][11] , \SB_CORRECT[14][11] , 
        \DB_DETECT[14][11] , \ACCESS_BUSY[14][12] , 
        \SB_CORRECT[14][12] , \DB_DETECT[14][12] , 
        \ACCESS_BUSY[14][13] , \SB_CORRECT[14][13] , 
        \DB_DETECT[14][13] , \ACCESS_BUSY[14][14] , 
        \SB_CORRECT[14][14] , \DB_DETECT[14][14] , 
        \ACCESS_BUSY[14][15] , \SB_CORRECT[14][15] , 
        \DB_DETECT[14][15] , \ACCESS_BUSY[14][16] , 
        \SB_CORRECT[14][16] , \DB_DETECT[14][16] , 
        \ACCESS_BUSY[14][17] , \SB_CORRECT[14][17] , 
        \DB_DETECT[14][17] , \ACCESS_BUSY[14][18] , 
        \SB_CORRECT[14][18] , \DB_DETECT[14][18] , 
        \ACCESS_BUSY[14][19] , \SB_CORRECT[14][19] , 
        \DB_DETECT[14][19] , \ACCESS_BUSY[15][0] , \SB_CORRECT[15][0] , 
        \DB_DETECT[15][0] , \ACCESS_BUSY[15][1] , \SB_CORRECT[15][1] , 
        \DB_DETECT[15][1] , \ACCESS_BUSY[15][2] , \SB_CORRECT[15][2] , 
        \DB_DETECT[15][2] , \ACCESS_BUSY[15][3] , \SB_CORRECT[15][3] , 
        \DB_DETECT[15][3] , \ACCESS_BUSY[15][4] , \SB_CORRECT[15][4] , 
        \DB_DETECT[15][4] , \ACCESS_BUSY[15][5] , \SB_CORRECT[15][5] , 
        \DB_DETECT[15][5] , \ACCESS_BUSY[15][6] , \SB_CORRECT[15][6] , 
        \DB_DETECT[15][6] , \ACCESS_BUSY[15][7] , \SB_CORRECT[15][7] , 
        \DB_DETECT[15][7] , \ACCESS_BUSY[15][8] , \SB_CORRECT[15][8] , 
        \DB_DETECT[15][8] , \ACCESS_BUSY[15][9] , \SB_CORRECT[15][9] , 
        \DB_DETECT[15][9] , \ACCESS_BUSY[15][10] , 
        \SB_CORRECT[15][10] , \DB_DETECT[15][10] , 
        \ACCESS_BUSY[15][11] , \SB_CORRECT[15][11] , 
        \DB_DETECT[15][11] , \ACCESS_BUSY[15][12] , 
        \SB_CORRECT[15][12] , \DB_DETECT[15][12] , 
        \ACCESS_BUSY[15][13] , \SB_CORRECT[15][13] , 
        \DB_DETECT[15][13] , \ACCESS_BUSY[15][14] , 
        \SB_CORRECT[15][14] , \DB_DETECT[15][14] , 
        \ACCESS_BUSY[15][15] , \SB_CORRECT[15][15] , 
        \DB_DETECT[15][15] , \ACCESS_BUSY[15][16] , 
        \SB_CORRECT[15][16] , \DB_DETECT[15][16] , 
        \ACCESS_BUSY[15][17] , \SB_CORRECT[15][17] , 
        \DB_DETECT[15][17] , \ACCESS_BUSY[15][18] , 
        \SB_CORRECT[15][18] , \DB_DETECT[15][18] , 
        \ACCESS_BUSY[15][19] , \SB_CORRECT[15][19] , 
        \DB_DETECT[15][19] , \ACCESS_BUSY[16][0] , \SB_CORRECT[16][0] , 
        \DB_DETECT[16][0] , \ACCESS_BUSY[16][1] , \SB_CORRECT[16][1] , 
        \DB_DETECT[16][1] , \ACCESS_BUSY[16][2] , \SB_CORRECT[16][2] , 
        \DB_DETECT[16][2] , \ACCESS_BUSY[16][3] , \SB_CORRECT[16][3] , 
        \DB_DETECT[16][3] , \ACCESS_BUSY[16][4] , \SB_CORRECT[16][4] , 
        \DB_DETECT[16][4] , \ACCESS_BUSY[16][5] , \SB_CORRECT[16][5] , 
        \DB_DETECT[16][5] , \ACCESS_BUSY[16][6] , \SB_CORRECT[16][6] , 
        \DB_DETECT[16][6] , \ACCESS_BUSY[16][7] , \SB_CORRECT[16][7] , 
        \DB_DETECT[16][7] , \ACCESS_BUSY[16][8] , \SB_CORRECT[16][8] , 
        \DB_DETECT[16][8] , \ACCESS_BUSY[16][9] , \SB_CORRECT[16][9] , 
        \DB_DETECT[16][9] , \ACCESS_BUSY[16][10] , 
        \SB_CORRECT[16][10] , \DB_DETECT[16][10] , 
        \ACCESS_BUSY[16][11] , \SB_CORRECT[16][11] , 
        \DB_DETECT[16][11] , \ACCESS_BUSY[16][12] , 
        \SB_CORRECT[16][12] , \DB_DETECT[16][12] , 
        \ACCESS_BUSY[16][13] , \SB_CORRECT[16][13] , 
        \DB_DETECT[16][13] , \ACCESS_BUSY[16][14] , 
        \SB_CORRECT[16][14] , \DB_DETECT[16][14] , 
        \ACCESS_BUSY[16][15] , \SB_CORRECT[16][15] , 
        \DB_DETECT[16][15] , \ACCESS_BUSY[16][16] , 
        \SB_CORRECT[16][16] , \DB_DETECT[16][16] , 
        \ACCESS_BUSY[16][17] , \SB_CORRECT[16][17] , 
        \DB_DETECT[16][17] , \ACCESS_BUSY[16][18] , 
        \SB_CORRECT[16][18] , \DB_DETECT[16][18] , 
        \ACCESS_BUSY[16][19] , \SB_CORRECT[16][19] , 
        \DB_DETECT[16][19] , \ACCESS_BUSY[17][0] , \SB_CORRECT[17][0] , 
        \DB_DETECT[17][0] , \ACCESS_BUSY[17][1] , \SB_CORRECT[17][1] , 
        \DB_DETECT[17][1] , \ACCESS_BUSY[17][2] , \SB_CORRECT[17][2] , 
        \DB_DETECT[17][2] , \ACCESS_BUSY[17][3] , \SB_CORRECT[17][3] , 
        \DB_DETECT[17][3] , \ACCESS_BUSY[17][4] , \SB_CORRECT[17][4] , 
        \DB_DETECT[17][4] , \ACCESS_BUSY[17][5] , \SB_CORRECT[17][5] , 
        \DB_DETECT[17][5] , \ACCESS_BUSY[17][6] , \SB_CORRECT[17][6] , 
        \DB_DETECT[17][6] , \ACCESS_BUSY[17][7] , \SB_CORRECT[17][7] , 
        \DB_DETECT[17][7] , \ACCESS_BUSY[17][8] , \SB_CORRECT[17][8] , 
        \DB_DETECT[17][8] , \ACCESS_BUSY[17][9] , \SB_CORRECT[17][9] , 
        \DB_DETECT[17][9] , \ACCESS_BUSY[17][10] , 
        \SB_CORRECT[17][10] , \DB_DETECT[17][10] , 
        \ACCESS_BUSY[17][11] , \SB_CORRECT[17][11] , 
        \DB_DETECT[17][11] , \ACCESS_BUSY[17][12] , 
        \SB_CORRECT[17][12] , \DB_DETECT[17][12] , 
        \ACCESS_BUSY[17][13] , \SB_CORRECT[17][13] , 
        \DB_DETECT[17][13] , \ACCESS_BUSY[17][14] , 
        \SB_CORRECT[17][14] , \DB_DETECT[17][14] , 
        \ACCESS_BUSY[17][15] , \SB_CORRECT[17][15] , 
        \DB_DETECT[17][15] , \ACCESS_BUSY[17][16] , 
        \SB_CORRECT[17][16] , \DB_DETECT[17][16] , 
        \ACCESS_BUSY[17][17] , \SB_CORRECT[17][17] , 
        \DB_DETECT[17][17] , \ACCESS_BUSY[17][18] , 
        \SB_CORRECT[17][18] , \DB_DETECT[17][18] , 
        \ACCESS_BUSY[17][19] , \SB_CORRECT[17][19] , 
        \DB_DETECT[17][19] , \ACCESS_BUSY[18][0] , \SB_CORRECT[18][0] , 
        \DB_DETECT[18][0] , \ACCESS_BUSY[18][1] , \SB_CORRECT[18][1] , 
        \DB_DETECT[18][1] , \ACCESS_BUSY[18][2] , \SB_CORRECT[18][2] , 
        \DB_DETECT[18][2] , \ACCESS_BUSY[18][3] , \SB_CORRECT[18][3] , 
        \DB_DETECT[18][3] , \ACCESS_BUSY[18][4] , \SB_CORRECT[18][4] , 
        \DB_DETECT[18][4] , \ACCESS_BUSY[18][5] , \SB_CORRECT[18][5] , 
        \DB_DETECT[18][5] , \ACCESS_BUSY[18][6] , \SB_CORRECT[18][6] , 
        \DB_DETECT[18][6] , \ACCESS_BUSY[18][7] , \SB_CORRECT[18][7] , 
        \DB_DETECT[18][7] , \ACCESS_BUSY[18][8] , \SB_CORRECT[18][8] , 
        \DB_DETECT[18][8] , \ACCESS_BUSY[18][9] , \SB_CORRECT[18][9] , 
        \DB_DETECT[18][9] , \ACCESS_BUSY[18][10] , 
        \SB_CORRECT[18][10] , \DB_DETECT[18][10] , 
        \ACCESS_BUSY[18][11] , \SB_CORRECT[18][11] , 
        \DB_DETECT[18][11] , \ACCESS_BUSY[18][12] , 
        \SB_CORRECT[18][12] , \DB_DETECT[18][12] , 
        \ACCESS_BUSY[18][13] , \SB_CORRECT[18][13] , 
        \DB_DETECT[18][13] , \ACCESS_BUSY[18][14] , 
        \SB_CORRECT[18][14] , \DB_DETECT[18][14] , 
        \ACCESS_BUSY[18][15] , \SB_CORRECT[18][15] , 
        \DB_DETECT[18][15] , \ACCESS_BUSY[18][16] , 
        \SB_CORRECT[18][16] , \DB_DETECT[18][16] , 
        \ACCESS_BUSY[18][17] , \SB_CORRECT[18][17] , 
        \DB_DETECT[18][17] , \ACCESS_BUSY[18][18] , 
        \SB_CORRECT[18][18] , \DB_DETECT[18][18] , 
        \ACCESS_BUSY[18][19] , \SB_CORRECT[18][19] , 
        \DB_DETECT[18][19] , \ACCESS_BUSY[19][0] , \SB_CORRECT[19][0] , 
        \DB_DETECT[19][0] , \ACCESS_BUSY[19][1] , \SB_CORRECT[19][1] , 
        \DB_DETECT[19][1] , \ACCESS_BUSY[19][2] , \SB_CORRECT[19][2] , 
        \DB_DETECT[19][2] , \ACCESS_BUSY[19][3] , \SB_CORRECT[19][3] , 
        \DB_DETECT[19][3] , \ACCESS_BUSY[19][4] , \SB_CORRECT[19][4] , 
        \DB_DETECT[19][4] , \ACCESS_BUSY[19][5] , \SB_CORRECT[19][5] , 
        \DB_DETECT[19][5] , \ACCESS_BUSY[19][6] , \SB_CORRECT[19][6] , 
        \DB_DETECT[19][6] , \ACCESS_BUSY[19][7] , \SB_CORRECT[19][7] , 
        \DB_DETECT[19][7] , \ACCESS_BUSY[19][8] , \SB_CORRECT[19][8] , 
        \DB_DETECT[19][8] , \ACCESS_BUSY[19][9] , \SB_CORRECT[19][9] , 
        \DB_DETECT[19][9] , \ACCESS_BUSY[19][10] , 
        \SB_CORRECT[19][10] , \DB_DETECT[19][10] , 
        \ACCESS_BUSY[19][11] , \SB_CORRECT[19][11] , 
        \DB_DETECT[19][11] , \ACCESS_BUSY[19][12] , 
        \SB_CORRECT[19][12] , \DB_DETECT[19][12] , 
        \ACCESS_BUSY[19][13] , \SB_CORRECT[19][13] , 
        \DB_DETECT[19][13] , \ACCESS_BUSY[19][14] , 
        \SB_CORRECT[19][14] , \DB_DETECT[19][14] , 
        \ACCESS_BUSY[19][15] , \SB_CORRECT[19][15] , 
        \DB_DETECT[19][15] , \ACCESS_BUSY[19][16] , 
        \SB_CORRECT[19][16] , \DB_DETECT[19][16] , 
        \ACCESS_BUSY[19][17] , \SB_CORRECT[19][17] , 
        \DB_DETECT[19][17] , \ACCESS_BUSY[19][18] , 
        \SB_CORRECT[19][18] , \DB_DETECT[19][18] , 
        \ACCESS_BUSY[19][19] , \SB_CORRECT[19][19] , 
        \DB_DETECT[19][19] , \ACCESS_BUSY[20][0] , \SB_CORRECT[20][0] , 
        \DB_DETECT[20][0] , \ACCESS_BUSY[20][1] , \SB_CORRECT[20][1] , 
        \DB_DETECT[20][1] , \ACCESS_BUSY[20][2] , \SB_CORRECT[20][2] , 
        \DB_DETECT[20][2] , \ACCESS_BUSY[20][3] , \SB_CORRECT[20][3] , 
        \DB_DETECT[20][3] , \ACCESS_BUSY[20][4] , \SB_CORRECT[20][4] , 
        \DB_DETECT[20][4] , \ACCESS_BUSY[20][5] , \SB_CORRECT[20][5] , 
        \DB_DETECT[20][5] , \ACCESS_BUSY[20][6] , \SB_CORRECT[20][6] , 
        \DB_DETECT[20][6] , \ACCESS_BUSY[20][7] , \SB_CORRECT[20][7] , 
        \DB_DETECT[20][7] , \ACCESS_BUSY[20][8] , \SB_CORRECT[20][8] , 
        \DB_DETECT[20][8] , \ACCESS_BUSY[20][9] , \SB_CORRECT[20][9] , 
        \DB_DETECT[20][9] , \ACCESS_BUSY[20][10] , 
        \SB_CORRECT[20][10] , \DB_DETECT[20][10] , 
        \ACCESS_BUSY[20][11] , \SB_CORRECT[20][11] , 
        \DB_DETECT[20][11] , \ACCESS_BUSY[20][12] , 
        \SB_CORRECT[20][12] , \DB_DETECT[20][12] , 
        \ACCESS_BUSY[20][13] , \SB_CORRECT[20][13] , 
        \DB_DETECT[20][13] , \ACCESS_BUSY[20][14] , 
        \SB_CORRECT[20][14] , \DB_DETECT[20][14] , 
        \ACCESS_BUSY[20][15] , \SB_CORRECT[20][15] , 
        \DB_DETECT[20][15] , \ACCESS_BUSY[20][16] , 
        \SB_CORRECT[20][16] , \DB_DETECT[20][16] , 
        \ACCESS_BUSY[20][17] , \SB_CORRECT[20][17] , 
        \DB_DETECT[20][17] , \ACCESS_BUSY[20][18] , 
        \SB_CORRECT[20][18] , \DB_DETECT[20][18] , 
        \ACCESS_BUSY[20][19] , \SB_CORRECT[20][19] , 
        \DB_DETECT[20][19] , \ACCESS_BUSY[21][0] , \SB_CORRECT[21][0] , 
        \DB_DETECT[21][0] , \ACCESS_BUSY[21][1] , \SB_CORRECT[21][1] , 
        \DB_DETECT[21][1] , \ACCESS_BUSY[21][2] , \SB_CORRECT[21][2] , 
        \DB_DETECT[21][2] , \ACCESS_BUSY[21][3] , \SB_CORRECT[21][3] , 
        \DB_DETECT[21][3] , \ACCESS_BUSY[21][4] , \SB_CORRECT[21][4] , 
        \DB_DETECT[21][4] , \ACCESS_BUSY[21][5] , \SB_CORRECT[21][5] , 
        \DB_DETECT[21][5] , \ACCESS_BUSY[21][6] , \SB_CORRECT[21][6] , 
        \DB_DETECT[21][6] , \ACCESS_BUSY[21][7] , \SB_CORRECT[21][7] , 
        \DB_DETECT[21][7] , \ACCESS_BUSY[21][8] , \SB_CORRECT[21][8] , 
        \DB_DETECT[21][8] , \ACCESS_BUSY[21][9] , \SB_CORRECT[21][9] , 
        \DB_DETECT[21][9] , \ACCESS_BUSY[21][10] , 
        \SB_CORRECT[21][10] , \DB_DETECT[21][10] , 
        \ACCESS_BUSY[21][11] , \SB_CORRECT[21][11] , 
        \DB_DETECT[21][11] , \ACCESS_BUSY[21][12] , 
        \SB_CORRECT[21][12] , \DB_DETECT[21][12] , 
        \ACCESS_BUSY[21][13] , \SB_CORRECT[21][13] , 
        \DB_DETECT[21][13] , \ACCESS_BUSY[21][14] , 
        \SB_CORRECT[21][14] , \DB_DETECT[21][14] , 
        \ACCESS_BUSY[21][15] , \SB_CORRECT[21][15] , 
        \DB_DETECT[21][15] , \ACCESS_BUSY[21][16] , 
        \SB_CORRECT[21][16] , \DB_DETECT[21][16] , 
        \ACCESS_BUSY[21][17] , \SB_CORRECT[21][17] , 
        \DB_DETECT[21][17] , \ACCESS_BUSY[21][18] , 
        \SB_CORRECT[21][18] , \DB_DETECT[21][18] , 
        \ACCESS_BUSY[21][19] , \SB_CORRECT[21][19] , 
        \DB_DETECT[21][19] , \ACCESS_BUSY[22][0] , \SB_CORRECT[22][0] , 
        \DB_DETECT[22][0] , \ACCESS_BUSY[22][1] , \SB_CORRECT[22][1] , 
        \DB_DETECT[22][1] , \ACCESS_BUSY[22][2] , \SB_CORRECT[22][2] , 
        \DB_DETECT[22][2] , \ACCESS_BUSY[22][3] , \SB_CORRECT[22][3] , 
        \DB_DETECT[22][3] , \ACCESS_BUSY[22][4] , \SB_CORRECT[22][4] , 
        \DB_DETECT[22][4] , \ACCESS_BUSY[22][5] , \SB_CORRECT[22][5] , 
        \DB_DETECT[22][5] , \ACCESS_BUSY[22][6] , \SB_CORRECT[22][6] , 
        \DB_DETECT[22][6] , \ACCESS_BUSY[22][7] , \SB_CORRECT[22][7] , 
        \DB_DETECT[22][7] , \ACCESS_BUSY[22][8] , \SB_CORRECT[22][8] , 
        \DB_DETECT[22][8] , \ACCESS_BUSY[22][9] , \SB_CORRECT[22][9] , 
        \DB_DETECT[22][9] , \ACCESS_BUSY[22][10] , 
        \SB_CORRECT[22][10] , \DB_DETECT[22][10] , 
        \ACCESS_BUSY[22][11] , \SB_CORRECT[22][11] , 
        \DB_DETECT[22][11] , \ACCESS_BUSY[22][12] , 
        \SB_CORRECT[22][12] , \DB_DETECT[22][12] , 
        \ACCESS_BUSY[22][13] , \SB_CORRECT[22][13] , 
        \DB_DETECT[22][13] , \ACCESS_BUSY[22][14] , 
        \SB_CORRECT[22][14] , \DB_DETECT[22][14] , 
        \ACCESS_BUSY[22][15] , \SB_CORRECT[22][15] , 
        \DB_DETECT[22][15] , \ACCESS_BUSY[22][16] , 
        \SB_CORRECT[22][16] , \DB_DETECT[22][16] , 
        \ACCESS_BUSY[22][17] , \SB_CORRECT[22][17] , 
        \DB_DETECT[22][17] , \ACCESS_BUSY[22][18] , 
        \SB_CORRECT[22][18] , \DB_DETECT[22][18] , 
        \ACCESS_BUSY[22][19] , \SB_CORRECT[22][19] , 
        \DB_DETECT[22][19] , \ACCESS_BUSY[23][0] , \SB_CORRECT[23][0] , 
        \DB_DETECT[23][0] , \ACCESS_BUSY[23][1] , \SB_CORRECT[23][1] , 
        \DB_DETECT[23][1] , \ACCESS_BUSY[23][2] , \SB_CORRECT[23][2] , 
        \DB_DETECT[23][2] , \ACCESS_BUSY[23][3] , \SB_CORRECT[23][3] , 
        \DB_DETECT[23][3] , \ACCESS_BUSY[23][4] , \SB_CORRECT[23][4] , 
        \DB_DETECT[23][4] , \ACCESS_BUSY[23][5] , \SB_CORRECT[23][5] , 
        \DB_DETECT[23][5] , \ACCESS_BUSY[23][6] , \SB_CORRECT[23][6] , 
        \DB_DETECT[23][6] , \ACCESS_BUSY[23][7] , \SB_CORRECT[23][7] , 
        \DB_DETECT[23][7] , \ACCESS_BUSY[23][8] , \SB_CORRECT[23][8] , 
        \DB_DETECT[23][8] , \ACCESS_BUSY[23][9] , \SB_CORRECT[23][9] , 
        \DB_DETECT[23][9] , \ACCESS_BUSY[23][10] , 
        \SB_CORRECT[23][10] , \DB_DETECT[23][10] , 
        \ACCESS_BUSY[23][11] , \SB_CORRECT[23][11] , 
        \DB_DETECT[23][11] , \ACCESS_BUSY[23][12] , 
        \SB_CORRECT[23][12] , \DB_DETECT[23][12] , 
        \ACCESS_BUSY[23][13] , \SB_CORRECT[23][13] , 
        \DB_DETECT[23][13] , \ACCESS_BUSY[23][14] , 
        \SB_CORRECT[23][14] , \DB_DETECT[23][14] , 
        \ACCESS_BUSY[23][15] , \SB_CORRECT[23][15] , 
        \DB_DETECT[23][15] , \ACCESS_BUSY[23][16] , 
        \SB_CORRECT[23][16] , \DB_DETECT[23][16] , 
        \ACCESS_BUSY[23][17] , \SB_CORRECT[23][17] , 
        \DB_DETECT[23][17] , \ACCESS_BUSY[23][18] , 
        \SB_CORRECT[23][18] , \DB_DETECT[23][18] , 
        \ACCESS_BUSY[23][19] , \SB_CORRECT[23][19] , 
        \DB_DETECT[23][19] , \ACCESS_BUSY[24][0] , \SB_CORRECT[24][0] , 
        \DB_DETECT[24][0] , \ACCESS_BUSY[24][1] , \SB_CORRECT[24][1] , 
        \DB_DETECT[24][1] , \ACCESS_BUSY[24][2] , \SB_CORRECT[24][2] , 
        \DB_DETECT[24][2] , \ACCESS_BUSY[24][3] , \SB_CORRECT[24][3] , 
        \DB_DETECT[24][3] , \ACCESS_BUSY[24][4] , \SB_CORRECT[24][4] , 
        \DB_DETECT[24][4] , \ACCESS_BUSY[24][5] , \SB_CORRECT[24][5] , 
        \DB_DETECT[24][5] , \ACCESS_BUSY[24][6] , \SB_CORRECT[24][6] , 
        \DB_DETECT[24][6] , \ACCESS_BUSY[24][7] , \SB_CORRECT[24][7] , 
        \DB_DETECT[24][7] , \ACCESS_BUSY[24][8] , \SB_CORRECT[24][8] , 
        \DB_DETECT[24][8] , \ACCESS_BUSY[24][9] , \SB_CORRECT[24][9] , 
        \DB_DETECT[24][9] , \ACCESS_BUSY[24][10] , 
        \SB_CORRECT[24][10] , \DB_DETECT[24][10] , 
        \ACCESS_BUSY[24][11] , \SB_CORRECT[24][11] , 
        \DB_DETECT[24][11] , \ACCESS_BUSY[24][12] , 
        \SB_CORRECT[24][12] , \DB_DETECT[24][12] , 
        \ACCESS_BUSY[24][13] , \SB_CORRECT[24][13] , 
        \DB_DETECT[24][13] , \ACCESS_BUSY[24][14] , 
        \SB_CORRECT[24][14] , \DB_DETECT[24][14] , 
        \ACCESS_BUSY[24][15] , \SB_CORRECT[24][15] , 
        \DB_DETECT[24][15] , \ACCESS_BUSY[24][16] , 
        \SB_CORRECT[24][16] , \DB_DETECT[24][16] , 
        \ACCESS_BUSY[24][17] , \SB_CORRECT[24][17] , 
        \DB_DETECT[24][17] , \ACCESS_BUSY[24][18] , 
        \SB_CORRECT[24][18] , \DB_DETECT[24][18] , 
        \ACCESS_BUSY[24][19] , \SB_CORRECT[24][19] , 
        \DB_DETECT[24][19] , \ACCESS_BUSY[25][0] , \SB_CORRECT[25][0] , 
        \DB_DETECT[25][0] , \ACCESS_BUSY[25][1] , \SB_CORRECT[25][1] , 
        \DB_DETECT[25][1] , \ACCESS_BUSY[25][2] , \SB_CORRECT[25][2] , 
        \DB_DETECT[25][2] , \ACCESS_BUSY[25][3] , \SB_CORRECT[25][3] , 
        \DB_DETECT[25][3] , \ACCESS_BUSY[25][4] , \SB_CORRECT[25][4] , 
        \DB_DETECT[25][4] , \ACCESS_BUSY[25][5] , \SB_CORRECT[25][5] , 
        \DB_DETECT[25][5] , \ACCESS_BUSY[25][6] , \SB_CORRECT[25][6] , 
        \DB_DETECT[25][6] , \ACCESS_BUSY[25][7] , \SB_CORRECT[25][7] , 
        \DB_DETECT[25][7] , \ACCESS_BUSY[25][8] , \SB_CORRECT[25][8] , 
        \DB_DETECT[25][8] , \ACCESS_BUSY[25][9] , \SB_CORRECT[25][9] , 
        \DB_DETECT[25][9] , \ACCESS_BUSY[25][10] , 
        \SB_CORRECT[25][10] , \DB_DETECT[25][10] , 
        \ACCESS_BUSY[25][11] , \SB_CORRECT[25][11] , 
        \DB_DETECT[25][11] , \ACCESS_BUSY[25][12] , 
        \SB_CORRECT[25][12] , \DB_DETECT[25][12] , 
        \ACCESS_BUSY[25][13] , \SB_CORRECT[25][13] , 
        \DB_DETECT[25][13] , \ACCESS_BUSY[25][14] , 
        \SB_CORRECT[25][14] , \DB_DETECT[25][14] , 
        \ACCESS_BUSY[25][15] , \SB_CORRECT[25][15] , 
        \DB_DETECT[25][15] , \ACCESS_BUSY[25][16] , 
        \SB_CORRECT[25][16] , \DB_DETECT[25][16] , 
        \ACCESS_BUSY[25][17] , \SB_CORRECT[25][17] , 
        \DB_DETECT[25][17] , \ACCESS_BUSY[25][18] , 
        \SB_CORRECT[25][18] , \DB_DETECT[25][18] , 
        \ACCESS_BUSY[25][19] , \SB_CORRECT[25][19] , 
        \DB_DETECT[25][19] , \ACCESS_BUSY[26][0] , \SB_CORRECT[26][0] , 
        \DB_DETECT[26][0] , \ACCESS_BUSY[26][1] , \SB_CORRECT[26][1] , 
        \DB_DETECT[26][1] , \ACCESS_BUSY[26][2] , \SB_CORRECT[26][2] , 
        \DB_DETECT[26][2] , \ACCESS_BUSY[26][3] , \SB_CORRECT[26][3] , 
        \DB_DETECT[26][3] , \ACCESS_BUSY[26][4] , \SB_CORRECT[26][4] , 
        \DB_DETECT[26][4] , \ACCESS_BUSY[26][5] , \SB_CORRECT[26][5] , 
        \DB_DETECT[26][5] , \ACCESS_BUSY[26][6] , \SB_CORRECT[26][6] , 
        \DB_DETECT[26][6] , \ACCESS_BUSY[26][7] , \SB_CORRECT[26][7] , 
        \DB_DETECT[26][7] , \ACCESS_BUSY[26][8] , \SB_CORRECT[26][8] , 
        \DB_DETECT[26][8] , \ACCESS_BUSY[26][9] , \SB_CORRECT[26][9] , 
        \DB_DETECT[26][9] , \ACCESS_BUSY[26][10] , 
        \SB_CORRECT[26][10] , \DB_DETECT[26][10] , 
        \ACCESS_BUSY[26][11] , \SB_CORRECT[26][11] , 
        \DB_DETECT[26][11] , \ACCESS_BUSY[26][12] , 
        \SB_CORRECT[26][12] , \DB_DETECT[26][12] , 
        \ACCESS_BUSY[26][13] , \SB_CORRECT[26][13] , 
        \DB_DETECT[26][13] , \ACCESS_BUSY[26][14] , 
        \SB_CORRECT[26][14] , \DB_DETECT[26][14] , 
        \ACCESS_BUSY[26][15] , \SB_CORRECT[26][15] , 
        \DB_DETECT[26][15] , \ACCESS_BUSY[26][16] , 
        \SB_CORRECT[26][16] , \DB_DETECT[26][16] , 
        \ACCESS_BUSY[26][17] , \SB_CORRECT[26][17] , 
        \DB_DETECT[26][17] , \ACCESS_BUSY[26][18] , 
        \SB_CORRECT[26][18] , \DB_DETECT[26][18] , 
        \ACCESS_BUSY[26][19] , \SB_CORRECT[26][19] , 
        \DB_DETECT[26][19] , \ACCESS_BUSY[27][0] , \SB_CORRECT[27][0] , 
        \DB_DETECT[27][0] , \ACCESS_BUSY[27][1] , \SB_CORRECT[27][1] , 
        \DB_DETECT[27][1] , \ACCESS_BUSY[27][2] , \SB_CORRECT[27][2] , 
        \DB_DETECT[27][2] , \ACCESS_BUSY[27][3] , \SB_CORRECT[27][3] , 
        \DB_DETECT[27][3] , \ACCESS_BUSY[27][4] , \SB_CORRECT[27][4] , 
        \DB_DETECT[27][4] , \ACCESS_BUSY[27][5] , \SB_CORRECT[27][5] , 
        \DB_DETECT[27][5] , \ACCESS_BUSY[27][6] , \SB_CORRECT[27][6] , 
        \DB_DETECT[27][6] , \ACCESS_BUSY[27][7] , \SB_CORRECT[27][7] , 
        \DB_DETECT[27][7] , \ACCESS_BUSY[27][8] , \SB_CORRECT[27][8] , 
        \DB_DETECT[27][8] , \ACCESS_BUSY[27][9] , \SB_CORRECT[27][9] , 
        \DB_DETECT[27][9] , \ACCESS_BUSY[27][10] , 
        \SB_CORRECT[27][10] , \DB_DETECT[27][10] , 
        \ACCESS_BUSY[27][11] , \SB_CORRECT[27][11] , 
        \DB_DETECT[27][11] , \ACCESS_BUSY[27][12] , 
        \SB_CORRECT[27][12] , \DB_DETECT[27][12] , 
        \ACCESS_BUSY[27][13] , \SB_CORRECT[27][13] , 
        \DB_DETECT[27][13] , \ACCESS_BUSY[27][14] , 
        \SB_CORRECT[27][14] , \DB_DETECT[27][14] , 
        \ACCESS_BUSY[27][15] , \SB_CORRECT[27][15] , 
        \DB_DETECT[27][15] , \ACCESS_BUSY[27][16] , 
        \SB_CORRECT[27][16] , \DB_DETECT[27][16] , 
        \ACCESS_BUSY[27][17] , \SB_CORRECT[27][17] , 
        \DB_DETECT[27][17] , \ACCESS_BUSY[27][18] , 
        \SB_CORRECT[27][18] , \DB_DETECT[27][18] , 
        \ACCESS_BUSY[27][19] , \SB_CORRECT[27][19] , 
        \DB_DETECT[27][19] , \ACCESS_BUSY[28][0] , \SB_CORRECT[28][0] , 
        \DB_DETECT[28][0] , \ACCESS_BUSY[28][1] , \SB_CORRECT[28][1] , 
        \DB_DETECT[28][1] , \ACCESS_BUSY[28][2] , \SB_CORRECT[28][2] , 
        \DB_DETECT[28][2] , \ACCESS_BUSY[28][3] , \SB_CORRECT[28][3] , 
        \DB_DETECT[28][3] , \ACCESS_BUSY[28][4] , \SB_CORRECT[28][4] , 
        \DB_DETECT[28][4] , \ACCESS_BUSY[28][5] , \SB_CORRECT[28][5] , 
        \DB_DETECT[28][5] , \ACCESS_BUSY[28][6] , \SB_CORRECT[28][6] , 
        \DB_DETECT[28][6] , \ACCESS_BUSY[28][7] , \SB_CORRECT[28][7] , 
        \DB_DETECT[28][7] , \ACCESS_BUSY[28][8] , \SB_CORRECT[28][8] , 
        \DB_DETECT[28][8] , \ACCESS_BUSY[28][9] , \SB_CORRECT[28][9] , 
        \DB_DETECT[28][9] , \ACCESS_BUSY[28][10] , 
        \SB_CORRECT[28][10] , \DB_DETECT[28][10] , 
        \ACCESS_BUSY[28][11] , \SB_CORRECT[28][11] , 
        \DB_DETECT[28][11] , \ACCESS_BUSY[28][12] , 
        \SB_CORRECT[28][12] , \DB_DETECT[28][12] , 
        \ACCESS_BUSY[28][13] , \SB_CORRECT[28][13] , 
        \DB_DETECT[28][13] , \ACCESS_BUSY[28][14] , 
        \SB_CORRECT[28][14] , \DB_DETECT[28][14] , 
        \ACCESS_BUSY[28][15] , \SB_CORRECT[28][15] , 
        \DB_DETECT[28][15] , \ACCESS_BUSY[28][16] , 
        \SB_CORRECT[28][16] , \DB_DETECT[28][16] , 
        \ACCESS_BUSY[28][17] , \SB_CORRECT[28][17] , 
        \DB_DETECT[28][17] , \ACCESS_BUSY[28][18] , 
        \SB_CORRECT[28][18] , \DB_DETECT[28][18] , 
        \ACCESS_BUSY[28][19] , \SB_CORRECT[28][19] , 
        \DB_DETECT[28][19] , \ACCESS_BUSY[29][0] , \SB_CORRECT[29][0] , 
        \DB_DETECT[29][0] , \ACCESS_BUSY[29][1] , \SB_CORRECT[29][1] , 
        \DB_DETECT[29][1] , \ACCESS_BUSY[29][2] , \SB_CORRECT[29][2] , 
        \DB_DETECT[29][2] , \ACCESS_BUSY[29][3] , \SB_CORRECT[29][3] , 
        \DB_DETECT[29][3] , \ACCESS_BUSY[29][4] , \SB_CORRECT[29][4] , 
        \DB_DETECT[29][4] , \ACCESS_BUSY[29][5] , \SB_CORRECT[29][5] , 
        \DB_DETECT[29][5] , \ACCESS_BUSY[29][6] , \SB_CORRECT[29][6] , 
        \DB_DETECT[29][6] , \ACCESS_BUSY[29][7] , \SB_CORRECT[29][7] , 
        \DB_DETECT[29][7] , \ACCESS_BUSY[29][8] , \SB_CORRECT[29][8] , 
        \DB_DETECT[29][8] , \ACCESS_BUSY[29][9] , \SB_CORRECT[29][9] , 
        \DB_DETECT[29][9] , \ACCESS_BUSY[29][10] , 
        \SB_CORRECT[29][10] , \DB_DETECT[29][10] , 
        \ACCESS_BUSY[29][11] , \SB_CORRECT[29][11] , 
        \DB_DETECT[29][11] , \ACCESS_BUSY[29][12] , 
        \SB_CORRECT[29][12] , \DB_DETECT[29][12] , 
        \ACCESS_BUSY[29][13] , \SB_CORRECT[29][13] , 
        \DB_DETECT[29][13] , \ACCESS_BUSY[29][14] , 
        \SB_CORRECT[29][14] , \DB_DETECT[29][14] , 
        \ACCESS_BUSY[29][15] , \SB_CORRECT[29][15] , 
        \DB_DETECT[29][15] , \ACCESS_BUSY[29][16] , 
        \SB_CORRECT[29][16] , \DB_DETECT[29][16] , 
        \ACCESS_BUSY[29][17] , \SB_CORRECT[29][17] , 
        \DB_DETECT[29][17] , \ACCESS_BUSY[29][18] , 
        \SB_CORRECT[29][18] , \DB_DETECT[29][18] , 
        \ACCESS_BUSY[29][19] , \SB_CORRECT[29][19] , 
        \DB_DETECT[29][19] , \ACCESS_BUSY[30][0] , \SB_CORRECT[30][0] , 
        \DB_DETECT[30][0] , \ACCESS_BUSY[30][1] , \SB_CORRECT[30][1] , 
        \DB_DETECT[30][1] , \ACCESS_BUSY[30][2] , \SB_CORRECT[30][2] , 
        \DB_DETECT[30][2] , \ACCESS_BUSY[30][3] , \SB_CORRECT[30][3] , 
        \DB_DETECT[30][3] , \ACCESS_BUSY[30][4] , \SB_CORRECT[30][4] , 
        \DB_DETECT[30][4] , \ACCESS_BUSY[30][5] , \SB_CORRECT[30][5] , 
        \DB_DETECT[30][5] , \ACCESS_BUSY[30][6] , \SB_CORRECT[30][6] , 
        \DB_DETECT[30][6] , \ACCESS_BUSY[30][7] , \SB_CORRECT[30][7] , 
        \DB_DETECT[30][7] , \ACCESS_BUSY[30][8] , \SB_CORRECT[30][8] , 
        \DB_DETECT[30][8] , \ACCESS_BUSY[30][9] , \SB_CORRECT[30][9] , 
        \DB_DETECT[30][9] , \ACCESS_BUSY[30][10] , 
        \SB_CORRECT[30][10] , \DB_DETECT[30][10] , 
        \ACCESS_BUSY[30][11] , \SB_CORRECT[30][11] , 
        \DB_DETECT[30][11] , \ACCESS_BUSY[30][12] , 
        \SB_CORRECT[30][12] , \DB_DETECT[30][12] , 
        \ACCESS_BUSY[30][13] , \SB_CORRECT[30][13] , 
        \DB_DETECT[30][13] , \ACCESS_BUSY[30][14] , 
        \SB_CORRECT[30][14] , \DB_DETECT[30][14] , 
        \ACCESS_BUSY[30][15] , \SB_CORRECT[30][15] , 
        \DB_DETECT[30][15] , \ACCESS_BUSY[30][16] , 
        \SB_CORRECT[30][16] , \DB_DETECT[30][16] , 
        \ACCESS_BUSY[30][17] , \SB_CORRECT[30][17] , 
        \DB_DETECT[30][17] , \ACCESS_BUSY[30][18] , 
        \SB_CORRECT[30][18] , \DB_DETECT[30][18] , 
        \ACCESS_BUSY[30][19] , \SB_CORRECT[30][19] , 
        \DB_DETECT[30][19] , \ACCESS_BUSY[31][0] , \SB_CORRECT[31][0] , 
        \DB_DETECT[31][0] , \ACCESS_BUSY[31][1] , \SB_CORRECT[31][1] , 
        \DB_DETECT[31][1] , \ACCESS_BUSY[31][2] , \SB_CORRECT[31][2] , 
        \DB_DETECT[31][2] , \ACCESS_BUSY[31][3] , \SB_CORRECT[31][3] , 
        \DB_DETECT[31][3] , \ACCESS_BUSY[31][4] , \SB_CORRECT[31][4] , 
        \DB_DETECT[31][4] , \ACCESS_BUSY[31][5] , \SB_CORRECT[31][5] , 
        \DB_DETECT[31][5] , \ACCESS_BUSY[31][6] , \SB_CORRECT[31][6] , 
        \DB_DETECT[31][6] , \ACCESS_BUSY[31][7] , \SB_CORRECT[31][7] , 
        \DB_DETECT[31][7] , \ACCESS_BUSY[31][8] , \SB_CORRECT[31][8] , 
        \DB_DETECT[31][8] , \ACCESS_BUSY[31][9] , \SB_CORRECT[31][9] , 
        \DB_DETECT[31][9] , \ACCESS_BUSY[31][10] , 
        \SB_CORRECT[31][10] , \DB_DETECT[31][10] , 
        \ACCESS_BUSY[31][11] , \SB_CORRECT[31][11] , 
        \DB_DETECT[31][11] , \ACCESS_BUSY[31][12] , 
        \SB_CORRECT[31][12] , \DB_DETECT[31][12] , 
        \ACCESS_BUSY[31][13] , \SB_CORRECT[31][13] , 
        \DB_DETECT[31][13] , \ACCESS_BUSY[31][14] , 
        \SB_CORRECT[31][14] , \DB_DETECT[31][14] , 
        \ACCESS_BUSY[31][15] , \SB_CORRECT[31][15] , 
        \DB_DETECT[31][15] , \ACCESS_BUSY[31][16] , 
        \SB_CORRECT[31][16] , \DB_DETECT[31][16] , 
        \ACCESS_BUSY[31][17] , \SB_CORRECT[31][17] , 
        \DB_DETECT[31][17] , \ACCESS_BUSY[31][18] , 
        \SB_CORRECT[31][18] , \DB_DETECT[31][18] , 
        \ACCESS_BUSY[31][19] , \SB_CORRECT[31][19] , 
        \DB_DETECT[31][19] , OR4_174_Y, OR4_214_Y, OR4_134_Y, 
        OR4_269_Y, OR4_47_Y, OR4_75_Y, OR4_190_Y, OR4_71_Y, OR4_235_Y, 
        OR2_21_Y, OR4_77_Y, OR4_244_Y, OR4_339_Y, OR4_12_Y, OR4_109_Y, 
        OR4_303_Y, OR4_81_Y, OR4_250_Y, OR4_195_Y, OR2_24_Y, OR4_212_Y, 
        OR4_130_Y, OR4_114_Y, OR4_106_Y, OR4_336_Y, OR4_268_Y, 
        OR4_258_Y, OR4_126_Y, OR4_53_Y, OR2_38_Y, OR4_41_Y, OR4_118_Y, 
        OR4_203_Y, OR4_279_Y, OR4_116_Y, OR4_315_Y, OR4_197_Y, 
        OR4_78_Y, OR4_182_Y, OR2_3_Y, OR4_153_Y, OR4_329_Y, OR4_56_Y, 
        OR4_99_Y, OR4_184_Y, OR4_19_Y, OR4_159_Y, OR4_335_Y, OR4_281_Y, 
        OR2_30_Y, OR4_301_Y, OR4_205_Y, OR4_191_Y, OR4_176_Y, OR4_54_Y, 
        OR4_357_Y, OR4_348_Y, OR4_200_Y, OR4_137_Y, OR2_1_Y, OR4_160_Y, 
        OR4_2_Y, OR4_63_Y, OR4_86_Y, OR4_340_Y, OR4_229_Y, OR4_248_Y, 
        OR4_318_Y, OR4_91_Y, OR2_33_Y, OR4_40_Y, OR4_211_Y, OR4_306_Y, 
        OR4_347_Y, OR4_76_Y, OR4_276_Y, OR4_45_Y, OR4_219_Y, OR4_161_Y, 
        OR2_36_Y, OR4_187_Y, OR4_98_Y, OR4_79_Y, OR4_68_Y, OR4_305_Y, 
        OR4_233_Y, OR4_227_Y, OR4_93_Y, OR4_21_Y, OR2_10_Y, OR4_256_Y, 
        OR4_245_Y, OR4_196_Y, OR4_29_Y, OR4_324_Y, OR4_169_Y, 
        OR4_247_Y, OR4_72_Y, OR4_100_Y, OR2_0_Y, OR4_246_Y, OR4_88_Y, 
        OR4_142_Y, OR4_162_Y, OR4_57_Y, OR4_317_Y, OR4_333_Y, OR4_31_Y, 
        OR4_164_Y, OR2_37_Y, CFG2_3_Y, CFG2_6_Y, CFG2_1_Y, CFG2_5_Y, 
        OR4_345_Y, OR4_330_Y, OR4_282_Y, OR4_124_Y, OR4_42_Y, 
        OR4_257_Y, OR4_332_Y, OR4_147_Y, OR4_172_Y, OR2_6_Y, OR4_312_Y, 
        OR4_129_Y, OR4_263_Y, OR4_156_Y, OR4_96_Y, OR4_302_Y, 
        OR4_319_Y, OR4_136_Y, OR4_349_Y, OR2_7_Y, OR4_27_Y, OR4_204_Y, 
        OR4_352_Y, OR4_242_Y, OR4_168_Y, OR4_18_Y, OR4_34_Y, OR4_218_Y, 
        OR4_64_Y, OR2_14_Y, OR4_89_Y, OR4_180_Y, OR4_151_Y, OR4_179_Y, 
        OR4_110_Y, OR4_221_Y, OR4_316_Y, OR4_123_Y, OR4_139_Y, OR2_9_Y, 
        OR4_0_Y, OR4_346_Y, OR4_356_Y, OR4_237_Y, OR4_127_Y, OR4_178_Y, 
        OR4_177_Y, OR4_241_Y, OR4_92_Y, OR2_15_Y, OR4_135_Y, OR4_331_Y, 
        OR4_28_Y, OR4_48_Y, OR4_307_Y, OR4_199_Y, OR4_217_Y, OR4_289_Y, 
        OR4_49_Y, OR2_2_Y, OR4_51_Y, OR4_343_Y, OR4_222_Y, OR4_298_Y, 
        OR4_157_Y, OR4_288_Y, OR4_252_Y, OR4_112_Y, OR4_50_Y, OR2_5_Y, 
        OR4_117_Y, OR4_26_Y, OR4_9_Y, OR4_304_Y, OR4_254_Y, OR4_16_Y, 
        OR4_166_Y, OR4_322_Y, OR4_189_Y, OR2_28_Y, OR4_225_Y, 
        OR4_213_Y, OR4_163_Y, OR4_7_Y, OR4_296_Y, OR4_140_Y, OR4_216_Y, 
        OR4_36_Y, OR4_62_Y, OR2_16_Y, OR4_83_Y, OR4_61_Y, OR4_70_Y, 
        OR4_321_Y, OR4_201_Y, OR4_267_Y, OR4_265_Y, OR4_323_Y, 
        OR4_165_Y, OR2_19_Y, OR4_193_Y, OR4_122_Y, OR4_95_Y, OR4_22_Y, 
        OR4_341_Y, OR4_107_Y, OR4_253_Y, OR4_38_Y, OR4_277_Y, OR2_32_Y, 
        OR4_285_Y, OR4_97_Y, OR4_230_Y, OR4_133_Y, OR4_59_Y, OR4_275_Y, 
        OR4_290_Y, OR4_115_Y, OR4_313_Y, OR2_22_Y, OR4_192_Y, 
        OR4_170_Y, OR4_243_Y, OR4_274_Y, OR4_231_Y, OR4_113_Y, 
        OR4_234_Y, OR4_104_Y, OR4_240_Y, OR2_23_Y, OR4_328_Y, 
        OR4_311_Y, OR4_320_Y, OR4_202_Y, OR4_94_Y, OR4_146_Y, 
        OR4_145_Y, OR4_207_Y, OR4_52_Y, OR2_29_Y, OR4_278_Y, OR4_66_Y, 
        OR4_121_Y, OR4_149_Y, OR4_35_Y, OR4_111_Y, OR4_39_Y, OR4_226_Y, 
        OR4_20_Y, OR2_31_Y, OR4_84_Y, OR4_3_Y, OR4_338_Y, OR4_280_Y, 
        OR4_223_Y, OR4_355_Y, OR4_138_Y, OR4_291_Y, OR4_155_Y, 
        OR2_39_Y, OR4_342_Y, OR4_210_Y, OR4_23_Y, OR4_185_Y, OR4_286_Y, 
        OR4_359_Y, OR4_30_Y, OR4_300_Y, OR4_309_Y, OR2_12_Y, OR4_206_Y, 
        OR4_325_Y, OR4_224_Y, OR4_167_Y, OR4_350_Y, OR4_44_Y, 
        OR4_261_Y, OR4_215_Y, OR4_101_Y, OR2_25_Y, OR4_294_Y, OR4_13_Y, 
        OR4_171_Y, OR4_33_Y, OR4_266_Y, OR4_186_Y, OR4_270_Y, OR4_73_Y, 
        OR4_67_Y, OR2_4_Y, OR4_58_Y, OR4_299_Y, OR4_119_Y, OR4_271_Y, 
        OR4_5_Y, OR4_80_Y, OR4_125_Y, OR4_17_Y, OR4_25_Y, OR2_17_Y, 
        OR4_344_Y, OR4_295_Y, OR4_132_Y, OR4_173_Y, OR4_228_Y, 
        OR4_150_Y, OR4_102_Y, OR4_120_Y, OR4_108_Y, OR2_13_Y, OR4_14_Y, 
        OR4_103_Y, OR4_259_Y, OR4_128_Y, OR4_354_Y, OR4_272_Y, 
        OR4_358_Y, OR4_148_Y, OR4_144_Y, OR2_11_Y, OR4_82_Y, OR4_251_Y, 
        OR4_11_Y, OR4_55_Y, OR4_43_Y, OR4_158_Y, OR4_90_Y, OR4_87_Y, 
        OR4_69_Y, OR2_8_Y, OR4_297_Y, OR4_337_Y, OR4_220_Y, OR4_293_Y, 
        OR4_287_Y, OR4_283_Y, OR4_255_Y, OR4_353_Y, OR4_46_Y, OR2_35_Y, 
        OR4_60_Y, OR4_15_Y, OR4_208_Y, OR4_260_Y, OR4_314_Y, OR4_239_Y, 
        OR4_175_Y, OR4_194_Y, OR4_183_Y, OR2_18_Y, OR4_308_Y, 
        OR4_181_Y, OR4_1_Y, OR4_152_Y, OR4_249_Y, OR4_327_Y, OR4_8_Y, 
        OR4_273_Y, OR4_284_Y, OR2_26_Y, OR4_262_Y, OR4_351_Y, 
        OR4_141_Y, OR4_10_Y, OR4_232_Y, OR4_154_Y, OR4_238_Y, OR4_37_Y, 
        OR4_32_Y, OR2_20_Y, CFG2_4_Y, CFG2_2_Y, CFG2_7_Y, CFG2_0_Y, 
        OR4_310_Y, OR4_264_Y, OR4_105_Y, OR4_143_Y, OR4_198_Y, 
        OR4_131_Y, OR4_65_Y, OR4_85_Y, OR4_74_Y, OR2_27_Y, OR4_292_Y, 
        OR4_334_Y, OR4_236_Y, OR4_188_Y, OR4_326_Y, OR4_4_Y, OR4_24_Y, 
        OR4_6_Y, OR4_209_Y, OR2_34_Y, VCC, GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C19 (.A_DOUT({nc0, 
        nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, nc10, nc11, nc12, 
        nc13, nc14, nc15, nc16, nc17, \R_DATA_TEMPR1[39] , 
        \R_DATA_TEMPR1[38] }), .B_DOUT({nc18, nc19, nc20, nc21, nc22, 
        nc23, nc24, nc25, nc26, nc27, nc28, nc29, nc30, nc31, nc32, 
        nc33, nc34, nc35, nc36, nc37}), .DB_DETECT(\DB_DETECT[1][19] ), 
        .SB_CORRECT(\SB_CORRECT[1][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_253 (.A(\R_DATA_TEMPR8[39] ), .B(\R_DATA_TEMPR9[39] ), .C(
        \R_DATA_TEMPR10[39] ), .D(\R_DATA_TEMPR11[39] ), .Y(OR4_253_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C16 (.A_DOUT({nc38, 
        nc39, nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, nc48, 
        nc49, nc50, nc51, nc52, nc53, nc54, nc55, \R_DATA_TEMPR23[33] , 
        \R_DATA_TEMPR23[32] }), .B_DOUT({nc56, nc57, nc58, nc59, nc60, 
        nc61, nc62, nc63, nc64, nc65, nc66, nc67, nc68, nc69, nc70, 
        nc71, nc72, nc73, nc74, nc75}), .DB_DETECT(\DB_DETECT[23][16] )
        , .SB_CORRECT(\SB_CORRECT[23][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C15 (.A_DOUT({nc76, 
        nc77, nc78, nc79, nc80, nc81, nc82, nc83, nc84, nc85, nc86, 
        nc87, nc88, nc89, nc90, nc91, nc92, nc93, \R_DATA_TEMPR3[31] , 
        \R_DATA_TEMPR3[30] }), .B_DOUT({nc94, nc95, nc96, nc97, nc98, 
        nc99, nc100, nc101, nc102, nc103, nc104, nc105, nc106, nc107, 
        nc108, nc109, nc110, nc111, nc112, nc113}), .DB_DETECT(
        \DB_DETECT[3][15] ), .SB_CORRECT(\SB_CORRECT[3][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C15 (.A_DOUT({nc114, 
        nc115, nc116, nc117, nc118, nc119, nc120, nc121, nc122, nc123, 
        nc124, nc125, nc126, nc127, nc128, nc129, nc130, nc131, 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR31[30] }), .B_DOUT({nc132, 
        nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, nc141, 
        nc142, nc143, nc144, nc145, nc146, nc147, nc148, nc149, nc150, 
        nc151}), .DB_DETECT(\DB_DETECT[31][15] ), .SB_CORRECT(
        \SB_CORRECT[31][15] ), .ACCESS_BUSY(\ACCESS_BUSY[31][15] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[7] , R_ADDR[14], R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[7] , W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_181 (.A(OR4_284_Y), .B(OR2_26_Y), .C(\R_DATA_TEMPR22[24] ), 
        .D(\R_DATA_TEMPR23[24] ), .Y(OR4_181_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C14 (.A_DOUT({nc152, 
        nc153, nc154, nc155, nc156, nc157, nc158, nc159, nc160, nc161, 
        nc162, nc163, nc164, nc165, nc166, nc167, nc168, nc169, 
        \R_DATA_TEMPR24[29] , \R_DATA_TEMPR24[28] }), .B_DOUT({nc170, 
        nc171, nc172, nc173, nc174, nc175, nc176, nc177, nc178, nc179, 
        nc180, nc181, nc182, nc183, nc184, nc185, nc186, nc187, nc188, 
        nc189}), .DB_DETECT(\DB_DETECT[24][14] ), .SB_CORRECT(
        \SB_CORRECT[24][14] ), .ACCESS_BUSY(\ACCESS_BUSY[24][14] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[6] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_106 (.A(\R_DATA_TEMPR28[13] ), .B(\R_DATA_TEMPR29[13] ), 
        .C(\R_DATA_TEMPR30[13] ), .D(\R_DATA_TEMPR31[13] ), .Y(
        OR4_106_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[2]  (.A(CFG2_7_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[2] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C14 (.A_DOUT({nc190, 
        nc191, nc192, nc193, nc194, nc195, nc196, nc197, nc198, nc199, 
        nc200, nc201, nc202, nc203, nc204, nc205, nc206, nc207, 
        \R_DATA_TEMPR6[29] , \R_DATA_TEMPR6[28] }), .B_DOUT({nc208, 
        nc209, nc210, nc211, nc212, nc213, nc214, nc215, nc216, nc217, 
        nc218, nc219, nc220, nc221, nc222, nc223, nc224, nc225, nc226, 
        nc227}), .DB_DETECT(\DB_DETECT[6][14] ), .SB_CORRECT(
        \SB_CORRECT[6][14] ), .ACCESS_BUSY(\ACCESS_BUSY[6][14] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[1] , R_ADDR[14], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[1] , W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_83 (.A(OR4_201_Y), .B(OR4_267_Y), .C(OR4_265_Y), .D(
        OR4_323_Y), .Y(OR4_83_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1 (.A_DOUT({nc228, 
        nc229, nc230, nc231, nc232, nc233, nc234, nc235, nc236, nc237, 
        nc238, nc239, nc240, nc241, nc242, nc243, nc244, nc245, 
        \R_DATA_TEMPR2[3] , \R_DATA_TEMPR2[2] }), .B_DOUT({nc246, 
        nc247, nc248, nc249, nc250, nc251, nc252, nc253, nc254, nc255, 
        nc256, nc257, nc258, nc259, nc260, nc261, nc262, nc263, nc264, 
        nc265}), .DB_DETECT(\DB_DETECT[2][1] ), .SB_CORRECT(
        \SB_CORRECT[2][1] ), .ACCESS_BUSY(\ACCESS_BUSY[2][1] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[0] , R_ADDR[14], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[0] , W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C15 (.A_DOUT({nc266, 
        nc267, nc268, nc269, nc270, nc271, nc272, nc273, nc274, nc275, 
        nc276, nc277, nc278, nc279, nc280, nc281, nc282, nc283, 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR23[30] }), .B_DOUT({nc284, 
        nc285, nc286, nc287, nc288, nc289, nc290, nc291, nc292, nc293, 
        nc294, nc295, nc296, nc297, nc298, nc299, nc300, nc301, nc302, 
        nc303}), .DB_DETECT(\DB_DETECT[23][15] ), .SB_CORRECT(
        \SB_CORRECT[23][15] ), .ACCESS_BUSY(\ACCESS_BUSY[23][15] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[5] , R_ADDR[14], R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[5] , W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_138 (.A(\R_DATA_TEMPR8[29] ), .B(\R_DATA_TEMPR9[29] ), .C(
        \R_DATA_TEMPR10[29] ), .D(\R_DATA_TEMPR11[29] ), .Y(OR4_138_Y));
    OR4 OR4_176 (.A(\R_DATA_TEMPR28[33] ), .B(\R_DATA_TEMPR29[33] ), 
        .C(\R_DATA_TEMPR30[33] ), .D(\R_DATA_TEMPR31[33] ), .Y(
        OR4_176_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C14 (.A_DOUT({nc304, 
        nc305, nc306, nc307, nc308, nc309, nc310, nc311, nc312, nc313, 
        nc314, nc315, nc316, nc317, nc318, nc319, nc320, nc321, 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR25[28] }), .B_DOUT({nc322, 
        nc323, nc324, nc325, nc326, nc327, nc328, nc329, nc330, nc331, 
        nc332, nc333, nc334, nc335, nc336, nc337, nc338, nc339, nc340, 
        nc341}), .DB_DETECT(\DB_DETECT[25][14] ), .SB_CORRECT(
        \SB_CORRECT[25][14] ), .ACCESS_BUSY(\ACCESS_BUSY[25][14] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[6] , \BLKY1[0] , R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[6] , \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C4 (.A_DOUT({nc342, 
        nc343, nc344, nc345, nc346, nc347, nc348, nc349, nc350, nc351, 
        nc352, nc353, nc354, nc355, nc356, nc357, nc358, nc359, 
        \R_DATA_TEMPR5[9] , \R_DATA_TEMPR5[8] }), .B_DOUT({nc360, 
        nc361, nc362, nc363, nc364, nc365, nc366, nc367, nc368, nc369, 
        nc370, nc371, nc372, nc373, nc374, nc375, nc376, nc377, nc378, 
        nc379}), .DB_DETECT(\DB_DETECT[5][4] ), .SB_CORRECT(
        \SB_CORRECT[5][4] ), .ACCESS_BUSY(\ACCESS_BUSY[5][4] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[1] , \BLKY1[0] , R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[1] , \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C12 (.A_DOUT({nc380, 
        nc381, nc382, nc383, nc384, nc385, nc386, nc387, nc388, nc389, 
        nc390, nc391, nc392, nc393, nc394, nc395, nc396, nc397, 
        \R_DATA_TEMPR12[25] , \R_DATA_TEMPR12[24] }), .B_DOUT({nc398, 
        nc399, nc400, nc401, nc402, nc403, nc404, nc405, nc406, nc407, 
        nc408, nc409, nc410, nc411, nc412, nc413, nc414, nc415, nc416, 
        nc417}), .DB_DETECT(\DB_DETECT[12][12] ), .SB_CORRECT(
        \SB_CORRECT[12][12] ), .ACCESS_BUSY(\ACCESS_BUSY[12][12] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C11 (.A_DOUT({nc418, 
        nc419, nc420, nc421, nc422, nc423, nc424, nc425, nc426, nc427, 
        nc428, nc429, nc430, nc431, nc432, nc433, nc434, nc435, 
        \R_DATA_TEMPR22[23] , \R_DATA_TEMPR22[22] }), .B_DOUT({nc436, 
        nc437, nc438, nc439, nc440, nc441, nc442, nc443, nc444, nc445, 
        nc446, nc447, nc448, nc449, nc450, nc451, nc452, nc453, nc454, 
        nc455}), .DB_DETECT(\DB_DETECT[22][11] ), .SB_CORRECT(
        \SB_CORRECT[22][11] ), .ACCESS_BUSY(\ACCESS_BUSY[22][11] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[5] , R_ADDR[14], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[5] , W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_308 (.A(OR4_249_Y), .B(OR4_327_Y), .C(OR4_8_Y), .D(
        OR4_273_Y), .Y(OR4_308_Y));
    OR4 OR4_317 (.A(\R_DATA_TEMPR4[36] ), .B(\R_DATA_TEMPR5[36] ), .C(
        \R_DATA_TEMPR6[36] ), .D(\R_DATA_TEMPR7[36] ), .Y(OR4_317_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C9 (.A_DOUT({nc456, 
        nc457, nc458, nc459, nc460, nc461, nc462, nc463, nc464, nc465, 
        nc466, nc467, nc468, nc469, nc470, nc471, nc472, nc473, 
        \R_DATA_TEMPR6[19] , \R_DATA_TEMPR6[18] }), .B_DOUT({nc474, 
        nc475, nc476, nc477, nc478, nc479, nc480, nc481, nc482, nc483, 
        nc484, nc485, nc486, nc487, nc488, nc489, nc490, nc491, nc492, 
        nc493}), .DB_DETECT(\DB_DETECT[6][9] ), .SB_CORRECT(
        \SB_CORRECT[6][9] ), .ACCESS_BUSY(\ACCESS_BUSY[6][9] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[1] , R_ADDR[14], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[1] , W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_110 (.A(\R_DATA_TEMPR0[3] ), .B(\R_DATA_TEMPR1[3] ), .C(
        \R_DATA_TEMPR2[3] ), .D(\R_DATA_TEMPR3[3] ), .Y(OR4_110_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C13 (.A_DOUT({nc494, 
        nc495, nc496, nc497, nc498, nc499, nc500, nc501, nc502, nc503, 
        nc504, nc505, nc506, nc507, nc508, nc509, nc510, nc511, 
        \R_DATA_TEMPR20[27] , \R_DATA_TEMPR20[26] }), .B_DOUT({nc512, 
        nc513, nc514, nc515, nc516, nc517, nc518, nc519, nc520, nc521, 
        nc522, nc523, nc524, nc525, nc526, nc527, nc528, nc529, nc530, 
        nc531}), .DB_DETECT(\DB_DETECT[20][13] ), .SB_CORRECT(
        \SB_CORRECT[20][13] ), .ACCESS_BUSY(\ACCESS_BUSY[20][13] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[5] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C1 (.A_DOUT({nc532, 
        nc533, nc534, nc535, nc536, nc537, nc538, nc539, nc540, nc541, 
        nc542, nc543, nc544, nc545, nc546, nc547, nc548, nc549, 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR30[2] }), .B_DOUT({nc550, 
        nc551, nc552, nc553, nc554, nc555, nc556, nc557, nc558, nc559, 
        nc560, nc561, nc562, nc563, nc564, nc565, nc566, nc567, nc568, 
        nc569}), .DB_DETECT(\DB_DETECT[30][1] ), .SB_CORRECT(
        \SB_CORRECT[30][1] ), .ACCESS_BUSY(\ACCESS_BUSY[30][1] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[7] , R_ADDR[14], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[7] , W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C17 (.A_DOUT({nc570, 
        nc571, nc572, nc573, nc574, nc575, nc576, nc577, nc578, nc579, 
        nc580, nc581, nc582, nc583, nc584, nc585, nc586, nc587, 
        \R_DATA_TEMPR2[35] , \R_DATA_TEMPR2[34] }), .B_DOUT({nc588, 
        nc589, nc590, nc591, nc592, nc593, nc594, nc595, nc596, nc597, 
        nc598, nc599, nc600, nc601, nc602, nc603, nc604, nc605, nc606, 
        nc607}), .DB_DETECT(\DB_DETECT[2][17] ), .SB_CORRECT(
        \SB_CORRECT[2][17] ), .ACCESS_BUSY(\ACCESS_BUSY[2][17] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[0] , R_ADDR[14], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[0] , W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C19 (.A_DOUT({nc608, 
        nc609, nc610, nc611, nc612, nc613, nc614, nc615, nc616, nc617, 
        nc618, nc619, nc620, nc621, nc622, nc623, nc624, nc625, 
        \R_DATA_TEMPR28[39] , \R_DATA_TEMPR28[38] }), .B_DOUT({nc626, 
        nc627, nc628, nc629, nc630, nc631, nc632, nc633, nc634, nc635, 
        nc636, nc637, nc638, nc639, nc640, nc641, nc642, nc643, nc644, 
        nc645}), .DB_DETECT(\DB_DETECT[28][19] ), .SB_CORRECT(
        \SB_CORRECT[28][19] ), .ACCESS_BUSY(\ACCESS_BUSY[28][19] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[7] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2 (.A(OR4_91_Y), .B(OR2_33_Y), .C(\R_DATA_TEMPR22[16] ), 
        .D(\R_DATA_TEMPR23[16] ), .Y(OR4_2_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1 (.A_DOUT({nc646, 
        nc647, nc648, nc649, nc650, nc651, nc652, nc653, nc654, nc655, 
        nc656, nc657, nc658, nc659, nc660, nc661, nc662, nc663, 
        \R_DATA_TEMPR7[3] , \R_DATA_TEMPR7[2] }), .B_DOUT({nc664, 
        nc665, nc666, nc667, nc668, nc669, nc670, nc671, nc672, nc673, 
        nc674, nc675, nc676, nc677, nc678, nc679, nc680, nc681, nc682, 
        nc683}), .DB_DETECT(\DB_DETECT[7][1] ), .SB_CORRECT(
        \SB_CORRECT[7][1] ), .ACCESS_BUSY(\ACCESS_BUSY[7][1] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[1] , R_ADDR[14], R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[1] , W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_329 (.A(OR4_281_Y), .B(OR2_30_Y), .C(\R_DATA_TEMPR22[37] ), 
        .D(\R_DATA_TEMPR23[37] ), .Y(OR4_329_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C5 (.A_DOUT({nc684, 
        nc685, nc686, nc687, nc688, nc689, nc690, nc691, nc692, nc693, 
        nc694, nc695, nc696, nc697, nc698, nc699, nc700, nc701, 
        \R_DATA_TEMPR16[11] , \R_DATA_TEMPR16[10] }), .B_DOUT({nc702, 
        nc703, nc704, nc705, nc706, nc707, nc708, nc709, nc710, nc711, 
        nc712, nc713, nc714, nc715, nc716, nc717, nc718, nc719, nc720, 
        nc721}), .DB_DETECT(\DB_DETECT[16][5] ), .SB_CORRECT(
        \SB_CORRECT[16][5] ), .ACCESS_BUSY(\ACCESS_BUSY[16][5] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[4] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C6 (.A_DOUT({nc722, 
        nc723, nc724, nc725, nc726, nc727, nc728, nc729, nc730, nc731, 
        nc732, nc733, nc734, nc735, nc736, nc737, nc738, nc739, 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR23[12] }), .B_DOUT({nc740, 
        nc741, nc742, nc743, nc744, nc745, nc746, nc747, nc748, nc749, 
        nc750, nc751, nc752, nc753, nc754, nc755, nc756, nc757, nc758, 
        nc759}), .DB_DETECT(\DB_DETECT[23][6] ), .SB_CORRECT(
        \SB_CORRECT[23][6] ), .ACCESS_BUSY(\ACCESS_BUSY[23][6] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[5] , R_ADDR[14], R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[5] , W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[29]  (.A(OR4_84_Y), .B(OR4_3_Y), .C(OR4_338_Y), .D(
        OR4_280_Y), .Y(R_DATA[29]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C4 (.A_DOUT({nc760, 
        nc761, nc762, nc763, nc764, nc765, nc766, nc767, nc768, nc769, 
        nc770, nc771, nc772, nc773, nc774, nc775, nc776, nc777, 
        \R_DATA_TEMPR1[9] , \R_DATA_TEMPR1[8] }), .B_DOUT({nc778, 
        nc779, nc780, nc781, nc782, nc783, nc784, nc785, nc786, nc787, 
        nc788, nc789, nc790, nc791, nc792, nc793, nc794, nc795, nc796, 
        nc797}), .DB_DETECT(\DB_DETECT[1][4] ), .SB_CORRECT(
        \SB_CORRECT[1][4] ), .ACCESS_BUSY(\ACCESS_BUSY[1][4] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[0] , \BLKY1[0] , R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[0] , \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C19 (.A_DOUT({nc798, 
        nc799, nc800, nc801, nc802, nc803, nc804, nc805, nc806, nc807, 
        nc808, nc809, nc810, nc811, nc812, nc813, nc814, nc815, 
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR8[38] }), .B_DOUT({nc816, 
        nc817, nc818, nc819, nc820, nc821, nc822, nc823, nc824, nc825, 
        nc826, nc827, nc828, nc829, nc830, nc831, nc832, nc833, nc834, 
        nc835}), .DB_DETECT(\DB_DETECT[8][19] ), .SB_CORRECT(
        \SB_CORRECT[8][19] ), .ACCESS_BUSY(\ACCESS_BUSY[8][19] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0 (.A_DOUT({nc836, 
        nc837, nc838, nc839, nc840, nc841, nc842, nc843, nc844, nc845, 
        nc846, nc847, nc848, nc849, nc850, nc851, nc852, nc853, 
        \R_DATA_TEMPR22[1] , \R_DATA_TEMPR22[0] }), .B_DOUT({nc854, 
        nc855, nc856, nc857, nc858, nc859, nc860, nc861, nc862, nc863, 
        nc864, nc865, nc866, nc867, nc868, nc869, nc870, nc871, nc872, 
        nc873}), .DB_DETECT(\DB_DETECT[22][0] ), .SB_CORRECT(
        \SB_CORRECT[22][0] ), .ACCESS_BUSY(\ACCESS_BUSY[22][0] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[5] , R_ADDR[14], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[5] , W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_48 (.A(\R_DATA_TEMPR28[26] ), .B(\R_DATA_TEMPR29[26] ), .C(
        \R_DATA_TEMPR30[26] ), .D(\R_DATA_TEMPR31[26] ), .Y(OR4_48_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C17 (.A_DOUT({nc874, 
        nc875, nc876, nc877, nc878, nc879, nc880, nc881, nc882, nc883, 
        nc884, nc885, nc886, nc887, nc888, nc889, nc890, nc891, 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR19[34] }), .B_DOUT({nc892, 
        nc893, nc894, nc895, nc896, nc897, nc898, nc899, nc900, nc901, 
        nc902, nc903, nc904, nc905, nc906, nc907, nc908, nc909, nc910, 
        nc911}), .DB_DETECT(\DB_DETECT[19][17] ), .SB_CORRECT(
        \SB_CORRECT[19][17] ), .ACCESS_BUSY(\ACCESS_BUSY[19][17] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[4] , R_ADDR[14], R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[4] , W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0 (.A_DOUT({nc912, 
        nc913, nc914, nc915, nc916, nc917, nc918, nc919, nc920, nc921, 
        nc922, nc923, nc924, nc925, nc926, nc927, nc928, nc929, 
        \R_DATA_TEMPR3[1] , \R_DATA_TEMPR3[0] }), .B_DOUT({nc930, 
        nc931, nc932, nc933, nc934, nc935, nc936, nc937, nc938, nc939, 
        nc940, nc941, nc942, nc943, nc944, nc945, nc946, nc947, nc948, 
        nc949}), .DB_DETECT(\DB_DETECT[3][0] ), .SB_CORRECT(
        \SB_CORRECT[3][0] ), .ACCESS_BUSY(\ACCESS_BUSY[3][0] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[0] , R_ADDR[14], R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[0] , W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_33 (.A(\R_DATA_TEMPR20[16] ), .B(\R_DATA_TEMPR21[16] ), .Y(
        OR2_33_Y));
    OR4 OR4_109 (.A(\R_DATA_TEMPR0[17] ), .B(\R_DATA_TEMPR1[17] ), .C(
        \R_DATA_TEMPR2[17] ), .D(\R_DATA_TEMPR3[17] ), .Y(OR4_109_Y));
    OR4 OR4_241 (.A(\R_DATA_TEMPR12[11] ), .B(\R_DATA_TEMPR13[11] ), 
        .C(\R_DATA_TEMPR14[11] ), .D(\R_DATA_TEMPR15[11] ), .Y(
        OR4_241_Y));
    OR2 OR2_15 (.A(\R_DATA_TEMPR20[11] ), .B(\R_DATA_TEMPR21[11] ), .Y(
        OR2_15_Y));
    OR4 OR4_81 (.A(\R_DATA_TEMPR8[17] ), .B(\R_DATA_TEMPR9[17] ), .C(
        \R_DATA_TEMPR10[17] ), .D(\R_DATA_TEMPR11[17] ), .Y(OR4_81_Y));
    OR4 OR4_118 (.A(OR4_182_Y), .B(OR2_3_Y), .C(\R_DATA_TEMPR22[9] ), 
        .D(\R_DATA_TEMPR23[9] ), .Y(OR4_118_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_206_Y), .B(OR4_325_Y), .C(OR4_224_Y), 
        .D(OR4_167_Y), .Y(R_DATA[7]));
    OR4 OR4_179 (.A(\R_DATA_TEMPR28[3] ), .B(\R_DATA_TEMPR29[3] ), .C(
        \R_DATA_TEMPR30[3] ), .D(\R_DATA_TEMPR31[3] ), .Y(OR4_179_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C5 (.A_DOUT({nc950, 
        nc951, nc952, nc953, nc954, nc955, nc956, nc957, nc958, nc959, 
        nc960, nc961, nc962, nc963, nc964, nc965, nc966, nc967, 
        \R_DATA_TEMPR28[11] , \R_DATA_TEMPR28[10] }), .B_DOUT({nc968, 
        nc969, nc970, nc971, nc972, nc973, nc974, nc975, nc976, nc977, 
        nc978, nc979, nc980, nc981, nc982, nc983, nc984, nc985, nc986, 
        nc987}), .DB_DETECT(\DB_DETECT[28][5] ), .SB_CORRECT(
        \SB_CORRECT[28][5] ), .ACCESS_BUSY(\ACCESS_BUSY[28][5] ), 
        .A_ADDR({R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], 
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({
        \BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, 
        GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], 
        W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({
        \BLKX2[7] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), 
        .B_WEN({GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C17 (.A_DOUT({nc988, 
        nc989, nc990, nc991, nc992, nc993, nc994, nc995, nc996, nc997, 
        nc998, nc999, nc1000, nc1001, nc1002, nc1003, nc1004, nc1005, 
        \R_DATA_TEMPR7[35] , \R_DATA_TEMPR7[34] }), .B_DOUT({nc1006, 
        nc1007, nc1008, nc1009, nc1010, nc1011, nc1012, nc1013, nc1014, 
        nc1015, nc1016, nc1017, nc1018, nc1019, nc1020, nc1021, nc1022, 
        nc1023, nc1024, nc1025}), .DB_DETECT(\DB_DETECT[7][17] ), 
        .SB_CORRECT(\SB_CORRECT[7][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C18 (.A_DOUT({
        nc1026, nc1027, nc1028, nc1029, nc1030, nc1031, nc1032, nc1033, 
        nc1034, nc1035, nc1036, nc1037, nc1038, nc1039, nc1040, nc1041, 
        nc1042, nc1043, \R_DATA_TEMPR28[37] , \R_DATA_TEMPR28[36] }), 
        .B_DOUT({nc1044, nc1045, nc1046, nc1047, nc1048, nc1049, 
        nc1050, nc1051, nc1052, nc1053, nc1054, nc1055, nc1056, nc1057, 
        nc1058, nc1059, nc1060, nc1061, nc1062, nc1063}), .DB_DETECT(
        \DB_DETECT[28][18] ), .SB_CORRECT(\SB_CORRECT[28][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C16 (.A_DOUT({
        nc1064, nc1065, nc1066, nc1067, nc1068, nc1069, nc1070, nc1071, 
        nc1072, nc1073, nc1074, nc1075, nc1076, nc1077, nc1078, nc1079, 
        nc1080, nc1081, \R_DATA_TEMPR20[33] , \R_DATA_TEMPR20[32] }), 
        .B_DOUT({nc1082, nc1083, nc1084, nc1085, nc1086, nc1087, 
        nc1088, nc1089, nc1090, nc1091, nc1092, nc1093, nc1094, nc1095, 
        nc1096, nc1097, nc1098, nc1099, nc1100, nc1101}), .DB_DETECT(
        \DB_DETECT[20][16] ), .SB_CORRECT(\SB_CORRECT[20][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C3 (.A_DOUT({nc1102, 
        nc1103, nc1104, nc1105, nc1106, nc1107, nc1108, nc1109, nc1110, 
        nc1111, nc1112, nc1113, nc1114, nc1115, nc1116, nc1117, nc1118, 
        nc1119, \R_DATA_TEMPR12[7] , \R_DATA_TEMPR12[6] }), .B_DOUT({
        nc1120, nc1121, nc1122, nc1123, nc1124, nc1125, nc1126, nc1127, 
        nc1128, nc1129, nc1130, nc1131, nc1132, nc1133, nc1134, nc1135, 
        nc1136, nc1137, nc1138, nc1139}), .DB_DETECT(
        \DB_DETECT[12][3] ), .SB_CORRECT(\SB_CORRECT[12][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1 (.A_DOUT({nc1140, 
        nc1141, nc1142, nc1143, nc1144, nc1145, nc1146, nc1147, nc1148, 
        nc1149, nc1150, nc1151, nc1152, nc1153, nc1154, nc1155, nc1156, 
        nc1157, \R_DATA_TEMPR5[3] , \R_DATA_TEMPR5[2] }), .B_DOUT({
        nc1158, nc1159, nc1160, nc1161, nc1162, nc1163, nc1164, nc1165, 
        nc1166, nc1167, nc1168, nc1169, nc1170, nc1171, nc1172, nc1173, 
        nc1174, nc1175, nc1176, nc1177}), .DB_DETECT(\DB_DETECT[5][1] )
        , .SB_CORRECT(\SB_CORRECT[5][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C14 (.A_DOUT({
        nc1178, nc1179, nc1180, nc1181, nc1182, nc1183, nc1184, nc1185, 
        nc1186, nc1187, nc1188, nc1189, nc1190, nc1191, nc1192, nc1193, 
        nc1194, nc1195, \R_DATA_TEMPR11[29] , \R_DATA_TEMPR11[28] }), 
        .B_DOUT({nc1196, nc1197, nc1198, nc1199, nc1200, nc1201, 
        nc1202, nc1203, nc1204, nc1205, nc1206, nc1207, nc1208, nc1209, 
        nc1210, nc1211, nc1212, nc1213, nc1214, nc1215}), .DB_DETECT(
        \DB_DETECT[11][14] ), .SB_CORRECT(\SB_CORRECT[11][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C13 (.A_DOUT({
        nc1216, nc1217, nc1218, nc1219, nc1220, nc1221, nc1222, nc1223, 
        nc1224, nc1225, nc1226, nc1227, nc1228, nc1229, nc1230, nc1231, 
        nc1232, nc1233, \R_DATA_TEMPR24[27] , \R_DATA_TEMPR24[26] }), 
        .B_DOUT({nc1234, nc1235, nc1236, nc1237, nc1238, nc1239, 
        nc1240, nc1241, nc1242, nc1243, nc1244, nc1245, nc1246, nc1247, 
        nc1248, nc1249, nc1250, nc1251, nc1252, nc1253}), .DB_DETECT(
        \DB_DETECT[24][13] ), .SB_CORRECT(\SB_CORRECT[24][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[4]  (.A(OR4_278_Y), .B(OR4_66_Y), .C(OR4_121_Y), 
        .D(OR4_149_Y), .Y(R_DATA[4]));
    OR4 OR4_135 (.A(OR4_307_Y), .B(OR4_199_Y), .C(OR4_217_Y), .D(
        OR4_289_Y), .Y(OR4_135_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C18 (.A_DOUT({nc1254, 
        nc1255, nc1256, nc1257, nc1258, nc1259, nc1260, nc1261, nc1262, 
        nc1263, nc1264, nc1265, nc1266, nc1267, nc1268, nc1269, nc1270, 
        nc1271, \R_DATA_TEMPR6[37] , \R_DATA_TEMPR6[36] }), .B_DOUT({
        nc1272, nc1273, nc1274, nc1275, nc1276, nc1277, nc1278, nc1279, 
        nc1280, nc1281, nc1282, nc1283, nc1284, nc1285, nc1286, nc1287, 
        nc1288, nc1289, nc1290, nc1291}), .DB_DETECT(
        \DB_DETECT[6][18] ), .SB_CORRECT(\SB_CORRECT[6][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C15 (.A_DOUT({
        nc1292, nc1293, nc1294, nc1295, nc1296, nc1297, nc1298, nc1299, 
        nc1300, nc1301, nc1302, nc1303, nc1304, nc1305, nc1306, nc1307, 
        nc1308, nc1309, \R_DATA_TEMPR20[31] , \R_DATA_TEMPR20[30] }), 
        .B_DOUT({nc1310, nc1311, nc1312, nc1313, nc1314, nc1315, 
        nc1316, nc1317, nc1318, nc1319, nc1320, nc1321, nc1322, nc1323, 
        nc1324, nc1325, nc1326, nc1327, nc1328, nc1329}), .DB_DETECT(
        \DB_DETECT[20][15] ), .SB_CORRECT(\SB_CORRECT[20][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_31 (.A(\R_DATA_TEMPR20[4] ), .B(\R_DATA_TEMPR21[4] ), .Y(
        OR2_31_Y));
    OR4 OR4_267 (.A(\R_DATA_TEMPR4[31] ), .B(\R_DATA_TEMPR5[31] ), .C(
        \R_DATA_TEMPR6[31] ), .D(\R_DATA_TEMPR7[31] ), .Y(OR4_267_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C13 (.A_DOUT({
        nc1330, nc1331, nc1332, nc1333, nc1334, nc1335, nc1336, nc1337, 
        nc1338, nc1339, nc1340, nc1341, nc1342, nc1343, nc1344, nc1345, 
        nc1346, nc1347, \R_DATA_TEMPR25[27] , \R_DATA_TEMPR25[26] }), 
        .B_DOUT({nc1348, nc1349, nc1350, nc1351, nc1352, nc1353, 
        nc1354, nc1355, nc1356, nc1357, nc1358, nc1359, nc1360, nc1361, 
        nc1362, nc1363, nc1364, nc1365, nc1366, nc1367}), .DB_DETECT(
        \DB_DETECT[25][13] ), .SB_CORRECT(\SB_CORRECT[25][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_167 (.A(\R_DATA_TEMPR28[7] ), .B(\R_DATA_TEMPR29[7] ), .C(
        \R_DATA_TEMPR30[7] ), .D(\R_DATA_TEMPR31[7] ), .Y(OR4_167_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C10 (.A_DOUT({nc1368, 
        nc1369, nc1370, nc1371, nc1372, nc1373, nc1374, nc1375, nc1376, 
        nc1377, nc1378, nc1379, nc1380, nc1381, nc1382, nc1383, nc1384, 
        nc1385, \R_DATA_TEMPR3[21] , \R_DATA_TEMPR3[20] }), .B_DOUT({
        nc1386, nc1387, nc1388, nc1389, nc1390, nc1391, nc1392, nc1393, 
        nc1394, nc1395, nc1396, nc1397, nc1398, nc1399, nc1400, nc1401, 
        nc1402, nc1403, nc1404, nc1405}), .DB_DETECT(
        \DB_DETECT[3][10] ), .SB_CORRECT(\SB_CORRECT[3][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C6 (.A_DOUT({nc1406, 
        nc1407, nc1408, nc1409, nc1410, nc1411, nc1412, nc1413, nc1414, 
        nc1415, nc1416, nc1417, nc1418, nc1419, nc1420, nc1421, nc1422, 
        nc1423, \R_DATA_TEMPR8[13] , \R_DATA_TEMPR8[12] }), .B_DOUT({
        nc1424, nc1425, nc1426, nc1427, nc1428, nc1429, nc1430, nc1431, 
        nc1432, nc1433, nc1434, nc1435, nc1436, nc1437, nc1438, nc1439, 
        nc1440, nc1441, nc1442, nc1443}), .DB_DETECT(\DB_DETECT[8][6] )
        , .SB_CORRECT(\SB_CORRECT[8][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C17 (.A_DOUT({nc1444, 
        nc1445, nc1446, nc1447, nc1448, nc1449, nc1450, nc1451, nc1452, 
        nc1453, nc1454, nc1455, nc1456, nc1457, nc1458, nc1459, nc1460, 
        nc1461, \R_DATA_TEMPR5[35] , \R_DATA_TEMPR5[34] }), .B_DOUT({
        nc1462, nc1463, nc1464, nc1465, nc1466, nc1467, nc1468, nc1469, 
        nc1470, nc1471, nc1472, nc1473, nc1474, nc1475, nc1476, nc1477, 
        nc1478, nc1479, nc1480, nc1481}), .DB_DETECT(
        \DB_DETECT[5][17] ), .SB_CORRECT(\SB_CORRECT[5][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C6 (.A_DOUT({nc1482, 
        nc1483, nc1484, nc1485, nc1486, nc1487, nc1488, nc1489, nc1490, 
        nc1491, nc1492, nc1493, nc1494, nc1495, nc1496, nc1497, nc1498, 
        nc1499, \R_DATA_TEMPR7[13] , \R_DATA_TEMPR7[12] }), .B_DOUT({
        nc1500, nc1501, nc1502, nc1503, nc1504, nc1505, nc1506, nc1507, 
        nc1508, nc1509, nc1510, nc1511, nc1512, nc1513, nc1514, nc1515, 
        nc1516, nc1517, nc1518, nc1519}), .DB_DETECT(\DB_DETECT[7][6] )
        , .SB_CORRECT(\SB_CORRECT[7][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_186 (.A(\R_DATA_TEMPR4[10] ), .B(\R_DATA_TEMPR5[10] ), .C(
        \R_DATA_TEMPR6[10] ), .D(\R_DATA_TEMPR7[10] ), .Y(OR4_186_Y));
    OR4 OR4_341 (.A(\R_DATA_TEMPR0[39] ), .B(\R_DATA_TEMPR1[39] ), .C(
        \R_DATA_TEMPR2[39] ), .D(\R_DATA_TEMPR3[39] ), .Y(OR4_341_Y));
    OR4 OR4_235 (.A(\R_DATA_TEMPR16[8] ), .B(\R_DATA_TEMPR17[8] ), .C(
        \R_DATA_TEMPR18[8] ), .D(\R_DATA_TEMPR19[8] ), .Y(OR4_235_Y));
    OR2 OR2_29 (.A(\R_DATA_TEMPR20[21] ), .B(\R_DATA_TEMPR21[21] ), .Y(
        OR2_29_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C5 (.A_DOUT({nc1520, 
        nc1521, nc1522, nc1523, nc1524, nc1525, nc1526, nc1527, nc1528, 
        nc1529, nc1530, nc1531, nc1532, nc1533, nc1534, nc1535, nc1536, 
        nc1537, \R_DATA_TEMPR11[11] , \R_DATA_TEMPR11[10] }), .B_DOUT({
        nc1538, nc1539, nc1540, nc1541, nc1542, nc1543, nc1544, nc1545, 
        nc1546, nc1547, nc1548, nc1549, nc1550, nc1551, nc1552, nc1553, 
        nc1554, nc1555, nc1556, nc1557}), .DB_DETECT(
        \DB_DETECT[11][5] ), .SB_CORRECT(\SB_CORRECT[11][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C15 (.A_DOUT({nc1558, 
        nc1559, nc1560, nc1561, nc1562, nc1563, nc1564, nc1565, nc1566, 
        nc1567, nc1568, nc1569, nc1570, nc1571, nc1572, nc1573, nc1574, 
        nc1575, \R_DATA_TEMPR0[31] , \R_DATA_TEMPR0[30] }), .B_DOUT({
        nc1576, nc1577, nc1578, nc1579, nc1580, nc1581, nc1582, nc1583, 
        nc1584, nc1585, nc1586, nc1587, nc1588, nc1589, nc1590, nc1591, 
        nc1592, nc1593, nc1594, nc1595}), .DB_DETECT(
        \DB_DETECT[0][15] ), .SB_CORRECT(\SB_CORRECT[0][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C5 (.A_DOUT({nc1596, 
        nc1597, nc1598, nc1599, nc1600, nc1601, nc1602, nc1603, nc1604, 
        nc1605, nc1606, nc1607, nc1608, nc1609, nc1610, nc1611, nc1612, 
        nc1613, \R_DATA_TEMPR14[11] , \R_DATA_TEMPR14[10] }), .B_DOUT({
        nc1614, nc1615, nc1616, nc1617, nc1618, nc1619, nc1620, nc1621, 
        nc1622, nc1623, nc1624, nc1625, nc1626, nc1627, nc1628, nc1629, 
        nc1630, nc1631, nc1632, nc1633}), .DB_DETECT(
        \DB_DETECT[14][5] ), .SB_CORRECT(\SB_CORRECT[14][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_264 (.A(OR4_74_Y), .B(OR2_27_Y), .C(\R_DATA_TEMPR22[28] ), 
        .D(\R_DATA_TEMPR23[28] ), .Y(OR4_264_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C18 (.A_DOUT({
        nc1634, nc1635, nc1636, nc1637, nc1638, nc1639, nc1640, nc1641, 
        nc1642, nc1643, nc1644, nc1645, nc1646, nc1647, nc1648, nc1649, 
        nc1650, nc1651, \R_DATA_TEMPR13[37] , \R_DATA_TEMPR13[36] }), 
        .B_DOUT({nc1652, nc1653, nc1654, nc1655, nc1656, nc1657, 
        nc1658, nc1659, nc1660, nc1661, nc1662, nc1663, nc1664, nc1665, 
        nc1666, nc1667, nc1668, nc1669, nc1670, nc1671}), .DB_DETECT(
        \DB_DETECT[13][18] ), .SB_CORRECT(\SB_CORRECT[13][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C9 (.A_DOUT({nc1672, 
        nc1673, nc1674, nc1675, nc1676, nc1677, nc1678, nc1679, nc1680, 
        nc1681, nc1682, nc1683, nc1684, nc1685, nc1686, nc1687, nc1688, 
        nc1689, \R_DATA_TEMPR5[19] , \R_DATA_TEMPR5[18] }), .B_DOUT({
        nc1690, nc1691, nc1692, nc1693, nc1694, nc1695, nc1696, nc1697, 
        nc1698, nc1699, nc1700, nc1701, nc1702, nc1703, nc1704, nc1705, 
        nc1706, nc1707, nc1708, nc1709}), .DB_DETECT(\DB_DETECT[5][9] )
        , .SB_CORRECT(\SB_CORRECT[5][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C8 (.A_DOUT({nc1710, 
        nc1711, nc1712, nc1713, nc1714, nc1715, nc1716, nc1717, nc1718, 
        nc1719, nc1720, nc1721, nc1722, nc1723, nc1724, nc1725, nc1726, 
        nc1727, \R_DATA_TEMPR12[17] , \R_DATA_TEMPR12[16] }), .B_DOUT({
        nc1728, nc1729, nc1730, nc1731, nc1732, nc1733, nc1734, nc1735, 
        nc1736, nc1737, nc1738, nc1739, nc1740, nc1741, nc1742, nc1743, 
        nc1744, nc1745, nc1746, nc1747}), .DB_DETECT(
        \DB_DETECT[12][8] ), .SB_CORRECT(\SB_CORRECT[12][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C12 (.A_DOUT({
        nc1748, nc1749, nc1750, nc1751, nc1752, nc1753, nc1754, nc1755, 
        nc1756, nc1757, nc1758, nc1759, nc1760, nc1761, nc1762, nc1763, 
        nc1764, nc1765, \R_DATA_TEMPR28[25] , \R_DATA_TEMPR28[24] }), 
        .B_DOUT({nc1766, nc1767, nc1768, nc1769, nc1770, nc1771, 
        nc1772, nc1773, nc1774, nc1775, nc1776, nc1777, nc1778, nc1779, 
        nc1780, nc1781, nc1782, nc1783, nc1784, nc1785}), .DB_DETECT(
        \DB_DETECT[28][12] ), .SB_CORRECT(\SB_CORRECT[28][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_293 (.A(\R_DATA_TEMPR28[0] ), .B(\R_DATA_TEMPR29[0] ), .C(
        \R_DATA_TEMPR30[0] ), .D(\R_DATA_TEMPR31[0] ), .Y(OR4_293_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C10 (.A_DOUT({
        nc1786, nc1787, nc1788, nc1789, nc1790, nc1791, nc1792, nc1793, 
        nc1794, nc1795, nc1796, nc1797, nc1798, nc1799, nc1800, nc1801, 
        nc1802, nc1803, \R_DATA_TEMPR28[21] , \R_DATA_TEMPR28[20] }), 
        .B_DOUT({nc1804, nc1805, nc1806, nc1807, nc1808, nc1809, 
        nc1810, nc1811, nc1812, nc1813, nc1814, nc1815, nc1816, nc1817, 
        nc1818, nc1819, nc1820, nc1821, nc1822, nc1823}), .DB_DETECT(
        \DB_DETECT[28][10] ), .SB_CORRECT(\SB_CORRECT[28][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C16 (.A_DOUT({
        nc1824, nc1825, nc1826, nc1827, nc1828, nc1829, nc1830, nc1831, 
        nc1832, nc1833, nc1834, nc1835, nc1836, nc1837, nc1838, nc1839, 
        nc1840, nc1841, \R_DATA_TEMPR24[33] , \R_DATA_TEMPR24[32] }), 
        .B_DOUT({nc1842, nc1843, nc1844, nc1845, nc1846, nc1847, 
        nc1848, nc1849, nc1850, nc1851, nc1852, nc1853, nc1854, nc1855, 
        nc1856, nc1857, nc1858, nc1859, nc1860, nc1861}), .DB_DETECT(
        \DB_DETECT[24][16] ), .SB_CORRECT(\SB_CORRECT[24][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C13 (.A_DOUT({nc1862, 
        nc1863, nc1864, nc1865, nc1866, nc1867, nc1868, nc1869, nc1870, 
        nc1871, nc1872, nc1873, nc1874, nc1875, nc1876, nc1877, nc1878, 
        nc1879, \R_DATA_TEMPR2[27] , \R_DATA_TEMPR2[26] }), .B_DOUT({
        nc1880, nc1881, nc1882, nc1883, nc1884, nc1885, nc1886, nc1887, 
        nc1888, nc1889, nc1890, nc1891, nc1892, nc1893, nc1894, nc1895, 
        nc1896, nc1897, nc1898, nc1899}), .DB_DETECT(
        \DB_DETECT[2][13] ), .SB_CORRECT(\SB_CORRECT[2][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_115 (.A(\R_DATA_TEMPR12[25] ), .B(\R_DATA_TEMPR13[25] ), 
        .C(\R_DATA_TEMPR14[25] ), .D(\R_DATA_TEMPR15[25] ), .Y(
        OR4_115_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C5 (.A_DOUT({nc1900, 
        nc1901, nc1902, nc1903, nc1904, nc1905, nc1906, nc1907, nc1908, 
        nc1909, nc1910, nc1911, nc1912, nc1913, nc1914, nc1915, nc1916, 
        nc1917, \R_DATA_TEMPR20[11] , \R_DATA_TEMPR20[10] }), .B_DOUT({
        nc1918, nc1919, nc1920, nc1921, nc1922, nc1923, nc1924, nc1925, 
        nc1926, nc1927, nc1928, nc1929, nc1930, nc1931, nc1932, nc1933, 
        nc1934, nc1935, nc1936, nc1937}), .DB_DETECT(
        \DB_DETECT[20][5] ), .SB_CORRECT(\SB_CORRECT[20][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_66 (.A(OR4_20_Y), .B(OR2_31_Y), .C(\R_DATA_TEMPR22[4] ), 
        .D(\R_DATA_TEMPR23[4] ), .Y(OR4_66_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C16 (.A_DOUT({
        nc1938, nc1939, nc1940, nc1941, nc1942, nc1943, nc1944, nc1945, 
        nc1946, nc1947, nc1948, nc1949, nc1950, nc1951, nc1952, nc1953, 
        nc1954, nc1955, \R_DATA_TEMPR25[33] , \R_DATA_TEMPR25[32] }), 
        .B_DOUT({nc1956, nc1957, nc1958, nc1959, nc1960, nc1961, 
        nc1962, nc1963, nc1964, nc1965, nc1966, nc1967, nc1968, nc1969, 
        nc1970, nc1971, nc1972, nc1973, nc1974, nc1975}), .DB_DETECT(
        \DB_DETECT[25][16] ), .SB_CORRECT(\SB_CORRECT[25][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h1) )  CFG2_4 (.A(W_ADDR[16]), .B(W_ADDR[15]), .Y(
        CFG2_4_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C15 (.A_DOUT({
        nc1976, nc1977, nc1978, nc1979, nc1980, nc1981, nc1982, nc1983, 
        nc1984, nc1985, nc1986, nc1987, nc1988, nc1989, nc1990, nc1991, 
        nc1992, nc1993, \R_DATA_TEMPR24[31] , \R_DATA_TEMPR24[30] }), 
        .B_DOUT({nc1994, nc1995, nc1996, nc1997, nc1998, nc1999, 
        nc2000, nc2001, nc2002, nc2003, nc2004, nc2005, nc2006, nc2007, 
        nc2008, nc2009, nc2010, nc2011, nc2012, nc2013}), .DB_DETECT(
        \DB_DETECT[24][15] ), .SB_CORRECT(\SB_CORRECT[24][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_238 (.A(\R_DATA_TEMPR8[20] ), .B(\R_DATA_TEMPR9[20] ), .C(
        \R_DATA_TEMPR10[20] ), .D(\R_DATA_TEMPR11[20] ), .Y(OR4_238_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C5 (.A_DOUT({nc2014, 
        nc2015, nc2016, nc2017, nc2018, nc2019, nc2020, nc2021, nc2022, 
        nc2023, nc2024, nc2025, nc2026, nc2027, nc2028, nc2029, nc2030, 
        nc2031, \R_DATA_TEMPR1[11] , \R_DATA_TEMPR1[10] }), .B_DOUT({
        nc2032, nc2033, nc2034, nc2035, nc2036, nc2037, nc2038, nc2039, 
        nc2040, nc2041, nc2042, nc2043, nc2044, nc2045, nc2046, nc2047, 
        nc2048, nc2049, nc2050, nc2051}), .DB_DETECT(\DB_DETECT[1][5] )
        , .SB_CORRECT(\SB_CORRECT[1][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C16 (.A_DOUT({
        nc2052, nc2053, nc2054, nc2055, nc2056, nc2057, nc2058, nc2059, 
        nc2060, nc2061, nc2062, nc2063, nc2064, nc2065, nc2066, nc2067, 
        nc2068, nc2069, \R_DATA_TEMPR18[33] , \R_DATA_TEMPR18[32] }), 
        .B_DOUT({nc2070, nc2071, nc2072, nc2073, nc2074, nc2075, 
        nc2076, nc2077, nc2078, nc2079, nc2080, nc2081, nc2082, nc2083, 
        nc2084, nc2085, nc2086, nc2087, nc2088, nc2089}), .DB_DETECT(
        \DB_DETECT[18][16] ), .SB_CORRECT(\SB_CORRECT[18][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_8 (.A(\R_DATA_TEMPR20[6] ), .B(\R_DATA_TEMPR21[6] ), .Y(
        OR2_8_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C7 (.A_DOUT({nc2090, 
        nc2091, nc2092, nc2093, nc2094, nc2095, nc2096, nc2097, nc2098, 
        nc2099, nc2100, nc2101, nc2102, nc2103, nc2104, nc2105, nc2106, 
        nc2107, \R_DATA_TEMPR5[15] , \R_DATA_TEMPR5[14] }), .B_DOUT({
        nc2108, nc2109, nc2110, nc2111, nc2112, nc2113, nc2114, nc2115, 
        nc2116, nc2117, nc2118, nc2119, nc2120, nc2121, nc2122, nc2123, 
        nc2124, nc2125, nc2126, nc2127}), .DB_DETECT(\DB_DETECT[5][7] )
        , .SB_CORRECT(\SB_CORRECT[5][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C9 (.A_DOUT({nc2128, 
        nc2129, nc2130, nc2131, nc2132, nc2133, nc2134, nc2135, nc2136, 
        nc2137, nc2138, nc2139, nc2140, nc2141, nc2142, nc2143, nc2144, 
        nc2145, \R_DATA_TEMPR26[19] , \R_DATA_TEMPR26[18] }), .B_DOUT({
        nc2146, nc2147, nc2148, nc2149, nc2150, nc2151, nc2152, nc2153, 
        nc2154, nc2155, nc2156, nc2157, nc2158, nc2159, nc2160, nc2161, 
        nc2162, nc2163, nc2164, nc2165}), .DB_DETECT(
        \DB_DETECT[26][9] ), .SB_CORRECT(\SB_CORRECT[26][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C7 (.A_DOUT({nc2166, 
        nc2167, nc2168, nc2169, nc2170, nc2171, nc2172, nc2173, nc2174, 
        nc2175, nc2176, nc2177, nc2178, nc2179, nc2180, nc2181, nc2182, 
        nc2183, \R_DATA_TEMPR29[15] , \R_DATA_TEMPR29[14] }), .B_DOUT({
        nc2184, nc2185, nc2186, nc2187, nc2188, nc2189, nc2190, nc2191, 
        nc2192, nc2193, nc2194, nc2195, nc2196, nc2197, nc2198, nc2199, 
        nc2200, nc2201, nc2202, nc2203}), .DB_DETECT(
        \DB_DETECT[29][7] ), .SB_CORRECT(\SB_CORRECT[29][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][7] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0 (.A_DOUT({nc2204, 
        nc2205, nc2206, nc2207, nc2208, nc2209, nc2210, nc2211, nc2212, 
        nc2213, nc2214, nc2215, nc2216, nc2217, nc2218, nc2219, nc2220, 
        nc2221, \R_DATA_TEMPR21[1] , \R_DATA_TEMPR21[0] }), .B_DOUT({
        nc2222, nc2223, nc2224, nc2225, nc2226, nc2227, nc2228, nc2229, 
        nc2230, nc2231, nc2232, nc2233, nc2234, nc2235, nc2236, nc2237, 
        nc2238, nc2239, nc2240, nc2241}), .DB_DETECT(
        \DB_DETECT[21][0] ), .SB_CORRECT(\SB_CORRECT[21][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_189 (.A(\R_DATA_TEMPR16[19] ), .B(\R_DATA_TEMPR17[19] ), 
        .C(\R_DATA_TEMPR18[19] ), .D(\R_DATA_TEMPR19[19] ), .Y(
        OR4_189_Y));
    OR4 OR4_0 (.A(OR4_127_Y), .B(OR4_178_Y), .C(OR4_177_Y), .D(
        OR4_241_Y), .Y(OR4_0_Y));
    OR4 OR4_207 (.A(\R_DATA_TEMPR12[21] ), .B(\R_DATA_TEMPR13[21] ), 
        .C(\R_DATA_TEMPR14[21] ), .D(\R_DATA_TEMPR15[21] ), .Y(
        OR4_207_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C15 (.A_DOUT({
        nc2242, nc2243, nc2244, nc2245, nc2246, nc2247, nc2248, nc2249, 
        nc2250, nc2251, nc2252, nc2253, nc2254, nc2255, nc2256, nc2257, 
        nc2258, nc2259, \R_DATA_TEMPR25[31] , \R_DATA_TEMPR25[30] }), 
        .B_DOUT({nc2260, nc2261, nc2262, nc2263, nc2264, nc2265, 
        nc2266, nc2267, nc2268, nc2269, nc2270, nc2271, nc2272, nc2273, 
        nc2274, nc2275, nc2276, nc2277, nc2278, nc2279}), .DB_DETECT(
        \DB_DETECT[25][15] ), .SB_CORRECT(\SB_CORRECT[25][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_215 (.A(\R_DATA_TEMPR12[7] ), .B(\R_DATA_TEMPR13[7] ), .C(
        \R_DATA_TEMPR14[7] ), .D(\R_DATA_TEMPR15[7] ), .Y(OR4_215_Y));
    OR4 OR4_107 (.A(\R_DATA_TEMPR4[39] ), .B(\R_DATA_TEMPR5[39] ), .C(
        \R_DATA_TEMPR6[39] ), .D(\R_DATA_TEMPR7[39] ), .Y(OR4_107_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C13 (.A_DOUT({nc2280, 
        nc2281, nc2282, nc2283, nc2284, nc2285, nc2286, nc2287, nc2288, 
        nc2289, nc2290, nc2291, nc2292, nc2293, nc2294, nc2295, nc2296, 
        nc2297, \R_DATA_TEMPR7[27] , \R_DATA_TEMPR7[26] }), .B_DOUT({
        nc2298, nc2299, nc2300, nc2301, nc2302, nc2303, nc2304, nc2305, 
        nc2306, nc2307, nc2308, nc2309, nc2310, nc2311, nc2312, nc2313, 
        nc2314, nc2315, nc2316, nc2317}), .DB_DETECT(
        \DB_DETECT[7][13] ), .SB_CORRECT(\SB_CORRECT[7][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_277 (.A(\R_DATA_TEMPR16[39] ), .B(\R_DATA_TEMPR17[39] ), 
        .C(\R_DATA_TEMPR18[39] ), .D(\R_DATA_TEMPR19[39] ), .Y(
        OR4_277_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C12 (.A_DOUT({
        nc2318, nc2319, nc2320, nc2321, nc2322, nc2323, nc2324, nc2325, 
        nc2326, nc2327, nc2328, nc2329, nc2330, nc2331, nc2332, nc2333, 
        nc2334, nc2335, \R_DATA_TEMPR19[25] , \R_DATA_TEMPR19[24] }), 
        .B_DOUT({nc2336, nc2337, nc2338, nc2339, nc2340, nc2341, 
        nc2342, nc2343, nc2344, nc2345, nc2346, nc2347, nc2348, nc2349, 
        nc2350, nc2351, nc2352, nc2353, nc2354, nc2355}), .DB_DETECT(
        \DB_DETECT[19][12] ), .SB_CORRECT(\SB_CORRECT[19][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C11 (.A_DOUT({
        nc2356, nc2357, nc2358, nc2359, nc2360, nc2361, nc2362, nc2363, 
        nc2364, nc2365, nc2366, nc2367, nc2368, nc2369, nc2370, nc2371, 
        nc2372, nc2373, \R_DATA_TEMPR29[23] , \R_DATA_TEMPR29[22] }), 
        .B_DOUT({nc2374, nc2375, nc2376, nc2377, nc2378, nc2379, 
        nc2380, nc2381, nc2382, nc2383, nc2384, nc2385, nc2386, nc2387, 
        nc2388, nc2389, nc2390, nc2391, nc2392, nc2393}), .DB_DETECT(
        \DB_DETECT[29][11] ), .SB_CORRECT(\SB_CORRECT[29][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C19 (.A_DOUT({
        nc2394, nc2395, nc2396, nc2397, nc2398, nc2399, nc2400, nc2401, 
        nc2402, nc2403, nc2404, nc2405, nc2406, nc2407, nc2408, nc2409, 
        nc2410, nc2411, \R_DATA_TEMPR21[39] , \R_DATA_TEMPR21[38] }), 
        .B_DOUT({nc2412, nc2413, nc2414, nc2415, nc2416, nc2417, 
        nc2418, nc2419, nc2420, nc2421, nc2422, nc2423, nc2424, nc2425, 
        nc2426, nc2427, nc2428, nc2429, nc2430, nc2431}), .DB_DETECT(
        \DB_DETECT[21][19] ), .SB_CORRECT(\SB_CORRECT[21][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_95 (.A(\R_DATA_TEMPR24[39] ), .B(\R_DATA_TEMPR25[39] ), .C(
        \R_DATA_TEMPR26[39] ), .D(\R_DATA_TEMPR27[39] ), .Y(OR4_95_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1 (.A_DOUT({nc2432, 
        nc2433, nc2434, nc2435, nc2436, nc2437, nc2438, nc2439, nc2440, 
        nc2441, nc2442, nc2443, nc2444, nc2445, nc2446, nc2447, nc2448, 
        nc2449, \R_DATA_TEMPR13[3] , \R_DATA_TEMPR13[2] }), .B_DOUT({
        nc2450, nc2451, nc2452, nc2453, nc2454, nc2455, nc2456, nc2457, 
        nc2458, nc2459, nc2460, nc2461, nc2462, nc2463, nc2464, nc2465, 
        nc2466, nc2467, nc2468, nc2469}), .DB_DETECT(
        \DB_DETECT[13][1] ), .SB_CORRECT(\SB_CORRECT[13][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_22 (.A(\R_DATA_TEMPR20[25] ), .B(\R_DATA_TEMPR21[25] ), .Y(
        OR2_22_Y));
    OR4 OR4_177 (.A(\R_DATA_TEMPR8[11] ), .B(\R_DATA_TEMPR9[11] ), .C(
        \R_DATA_TEMPR10[11] ), .D(\R_DATA_TEMPR11[11] ), .Y(OR4_177_Y));
    OR4 \OR4_R_DATA[34]  (.A(OR4_58_Y), .B(OR4_299_Y), .C(OR4_119_Y), 
        .D(OR4_271_Y), .Y(R_DATA[34]));
    OR4 OR4_349 (.A(\R_DATA_TEMPR16[15] ), .B(\R_DATA_TEMPR17[15] ), 
        .C(\R_DATA_TEMPR18[15] ), .D(\R_DATA_TEMPR19[15] ), .Y(
        OR4_349_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C3 (.A_DOUT({nc2470, 
        nc2471, nc2472, nc2473, nc2474, nc2475, nc2476, nc2477, nc2478, 
        nc2479, nc2480, nc2481, nc2482, nc2483, nc2484, nc2485, nc2486, 
        nc2487, \R_DATA_TEMPR27[7] , \R_DATA_TEMPR27[6] }), .B_DOUT({
        nc2488, nc2489, nc2490, nc2491, nc2492, nc2493, nc2494, nc2495, 
        nc2496, nc2497, nc2498, nc2499, nc2500, nc2501, nc2502, nc2503, 
        nc2504, nc2505, nc2506, nc2507}), .DB_DETECT(
        \DB_DETECT[27][3] ), .SB_CORRECT(\SB_CORRECT[27][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_223 (.A(\R_DATA_TEMPR0[29] ), .B(\R_DATA_TEMPR1[29] ), .C(
        \R_DATA_TEMPR2[29] ), .D(\R_DATA_TEMPR3[29] ), .Y(OR4_223_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C19 (.A_DOUT({
        nc2508, nc2509, nc2510, nc2511, nc2512, nc2513, nc2514, nc2515, 
        nc2516, nc2517, nc2518, nc2519, nc2520, nc2521, nc2522, nc2523, 
        nc2524, nc2525, \R_DATA_TEMPR16[39] , \R_DATA_TEMPR16[38] }), 
        .B_DOUT({nc2526, nc2527, nc2528, nc2529, nc2530, nc2531, 
        nc2532, nc2533, nc2534, nc2535, nc2536, nc2537, nc2538, nc2539, 
        nc2540, nc2541, nc2542, nc2543, nc2544, nc2545}), .DB_DETECT(
        \DB_DETECT[16][19] ), .SB_CORRECT(\SB_CORRECT[16][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0 (.A_DOUT({nc2546, 
        nc2547, nc2548, nc2549, nc2550, nc2551, nc2552, nc2553, nc2554, 
        nc2555, nc2556, nc2557, nc2558, nc2559, nc2560, nc2561, nc2562, 
        nc2563, \R_DATA_TEMPR17[1] , \R_DATA_TEMPR17[0] }), .B_DOUT({
        nc2564, nc2565, nc2566, nc2567, nc2568, nc2569, nc2570, nc2571, 
        nc2572, nc2573, nc2574, nc2575, nc2576, nc2577, nc2578, nc2579, 
        nc2580, nc2581, nc2582, nc2583}), .DB_DETECT(
        \DB_DETECT[17][0] ), .SB_CORRECT(\SB_CORRECT[17][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_354 (.A(\R_DATA_TEMPR0[30] ), .B(\R_DATA_TEMPR1[30] ), .C(
        \R_DATA_TEMPR2[30] ), .D(\R_DATA_TEMPR3[30] ), .Y(OR4_354_Y));
    OR4 OR4_204 (.A(OR4_64_Y), .B(OR2_14_Y), .C(\R_DATA_TEMPR22[35] ), 
        .D(\R_DATA_TEMPR23[35] ), .Y(OR4_204_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C7 (.A_DOUT({nc2584, 
        nc2585, nc2586, nc2587, nc2588, nc2589, nc2590, nc2591, nc2592, 
        nc2593, nc2594, nc2595, nc2596, nc2597, nc2598, nc2599, nc2600, 
        nc2601, \R_DATA_TEMPR13[15] , \R_DATA_TEMPR13[14] }), .B_DOUT({
        nc2602, nc2603, nc2604, nc2605, nc2606, nc2607, nc2608, nc2609, 
        nc2610, nc2611, nc2612, nc2613, nc2614, nc2615, nc2616, nc2617, 
        nc2618, nc2619, nc2620, nc2621}), .DB_DETECT(
        \DB_DETECT[13][7] ), .SB_CORRECT(\SB_CORRECT[13][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][7] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_19 (.A(\R_DATA_TEMPR20[31] ), .B(\R_DATA_TEMPR21[31] ), .Y(
        OR2_19_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C2 (.A_DOUT({nc2622, 
        nc2623, nc2624, nc2625, nc2626, nc2627, nc2628, nc2629, nc2630, 
        nc2631, nc2632, nc2633, nc2634, nc2635, nc2636, nc2637, nc2638, 
        nc2639, \R_DATA_TEMPR1[5] , \R_DATA_TEMPR1[4] }), .B_DOUT({
        nc2640, nc2641, nc2642, nc2643, nc2644, nc2645, nc2646, nc2647, 
        nc2648, nc2649, nc2650, nc2651, nc2652, nc2653, nc2654, nc2655, 
        nc2656, nc2657, nc2658, nc2659}), .DB_DETECT(\DB_DETECT[1][2] )
        , .SB_CORRECT(\SB_CORRECT[1][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C7 (.A_DOUT({nc2660, 
        nc2661, nc2662, nc2663, nc2664, nc2665, nc2666, nc2667, nc2668, 
        nc2669, nc2670, nc2671, nc2672, nc2673, nc2674, nc2675, nc2676, 
        nc2677, \R_DATA_TEMPR8[15] , \R_DATA_TEMPR8[14] }), .B_DOUT({
        nc2678, nc2679, nc2680, nc2681, nc2682, nc2683, nc2684, nc2685, 
        nc2686, nc2687, nc2688, nc2689, nc2690, nc2691, nc2692, nc2693, 
        nc2694, nc2695, nc2696, nc2697}), .DB_DETECT(\DB_DETECT[8][7] )
        , .SB_CORRECT(\SB_CORRECT[8][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_274 (.A(\R_DATA_TEMPR28[2] ), .B(\R_DATA_TEMPR29[2] ), .C(
        \R_DATA_TEMPR30[2] ), .D(\R_DATA_TEMPR31[2] ), .Y(OR4_274_Y));
    OR4 OR4_151 (.A(\R_DATA_TEMPR24[3] ), .B(\R_DATA_TEMPR25[3] ), .C(
        \R_DATA_TEMPR26[3] ), .D(\R_DATA_TEMPR27[3] ), .Y(OR4_151_Y));
    OR4 OR4_218 (.A(\R_DATA_TEMPR12[35] ), .B(\R_DATA_TEMPR13[35] ), 
        .C(\R_DATA_TEMPR14[35] ), .D(\R_DATA_TEMPR15[35] ), .Y(
        OR4_218_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_225_Y), .B(OR4_213_Y), .C(OR4_163_Y), 
        .D(OR4_7_Y), .Y(R_DATA[22]));
    OR4 OR4_60 (.A(OR4_314_Y), .B(OR4_239_Y), .C(OR4_175_Y), .D(
        OR4_194_Y), .Y(OR4_60_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C13 (.A_DOUT({
        nc2698, nc2699, nc2700, nc2701, nc2702, nc2703, nc2704, nc2705, 
        nc2706, nc2707, nc2708, nc2709, nc2710, nc2711, nc2712, nc2713, 
        nc2714, nc2715, \R_DATA_TEMPR18[27] , \R_DATA_TEMPR18[26] }), 
        .B_DOUT({nc2716, nc2717, nc2718, nc2719, nc2720, nc2721, 
        nc2722, nc2723, nc2724, nc2725, nc2726, nc2727, nc2728, nc2729, 
        nc2730, nc2731, nc2732, nc2733, nc2734, nc2735}), .DB_DETECT(
        \DB_DETECT[18][13] ), .SB_CORRECT(\SB_CORRECT[18][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C18 (.A_DOUT({
        nc2736, nc2737, nc2738, nc2739, nc2740, nc2741, nc2742, nc2743, 
        nc2744, nc2745, nc2746, nc2747, nc2748, nc2749, nc2750, nc2751, 
        nc2752, nc2753, \R_DATA_TEMPR10[37] , \R_DATA_TEMPR10[36] }), 
        .B_DOUT({nc2754, nc2755, nc2756, nc2757, nc2758, nc2759, 
        nc2760, nc2761, nc2762, nc2763, nc2764, nc2765, nc2766, nc2767, 
        nc2768, nc2769, nc2770, nc2771, nc2772, nc2773}), .DB_DETECT(
        \DB_DETECT[10][18] ), .SB_CORRECT(\SB_CORRECT[10][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C4 (.A_DOUT({nc2774, 
        nc2775, nc2776, nc2777, nc2778, nc2779, nc2780, nc2781, nc2782, 
        nc2783, nc2784, nc2785, nc2786, nc2787, nc2788, nc2789, nc2790, 
        nc2791, \R_DATA_TEMPR11[9] , \R_DATA_TEMPR11[8] }), .B_DOUT({
        nc2792, nc2793, nc2794, nc2795, nc2796, nc2797, nc2798, nc2799, 
        nc2800, nc2801, nc2802, nc2803, nc2804, nc2805, nc2806, nc2807, 
        nc2808, nc2809, nc2810, nc2811}), .DB_DETECT(
        \DB_DETECT[11][4] ), .SB_CORRECT(\SB_CORRECT[11][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C13 (.A_DOUT({nc2812, 
        nc2813, nc2814, nc2815, nc2816, nc2817, nc2818, nc2819, nc2820, 
        nc2821, nc2822, nc2823, nc2824, nc2825, nc2826, nc2827, nc2828, 
        nc2829, \R_DATA_TEMPR5[27] , \R_DATA_TEMPR5[26] }), .B_DOUT({
        nc2830, nc2831, nc2832, nc2833, nc2834, nc2835, nc2836, nc2837, 
        nc2838, nc2839, nc2840, nc2841, nc2842, nc2843, nc2844, nc2845, 
        nc2846, nc2847, nc2848, nc2849}), .DB_DETECT(
        \DB_DETECT[5][13] ), .SB_CORRECT(\SB_CORRECT[5][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C18 (.A_DOUT({
        nc2850, nc2851, nc2852, nc2853, nc2854, nc2855, nc2856, nc2857, 
        nc2858, nc2859, nc2860, nc2861, nc2862, nc2863, nc2864, nc2865, 
        nc2866, nc2867, \R_DATA_TEMPR21[37] , \R_DATA_TEMPR21[36] }), 
        .B_DOUT({nc2868, nc2869, nc2870, nc2871, nc2872, nc2873, 
        nc2874, nc2875, nc2876, nc2877, nc2878, nc2879, nc2880, nc2881, 
        nc2882, nc2883, nc2884, nc2885, nc2886, nc2887}), .DB_DETECT(
        \DB_DETECT[21][18] ), .SB_CORRECT(\SB_CORRECT[21][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_67 (.A(\R_DATA_TEMPR16[10] ), .B(\R_DATA_TEMPR17[10] ), .C(
        \R_DATA_TEMPR18[10] ), .D(\R_DATA_TEMPR19[10] ), .Y(OR4_67_Y));
    OR4 OR4_305 (.A(\R_DATA_TEMPR0[23] ), .B(\R_DATA_TEMPR1[23] ), .C(
        \R_DATA_TEMPR2[23] ), .D(\R_DATA_TEMPR3[23] ), .Y(OR4_305_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1 (.A_DOUT({nc2888, 
        nc2889, nc2890, nc2891, nc2892, nc2893, nc2894, nc2895, nc2896, 
        nc2897, nc2898, nc2899, nc2900, nc2901, nc2902, nc2903, nc2904, 
        nc2905, \R_DATA_TEMPR1[3] , \R_DATA_TEMPR1[2] }), .B_DOUT({
        nc2906, nc2907, nc2908, nc2909, nc2910, nc2911, nc2912, nc2913, 
        nc2914, nc2915, nc2916, nc2917, nc2918, nc2919, nc2920, nc2921, 
        nc2922, nc2923, nc2924, nc2925}), .DB_DETECT(\DB_DETECT[1][1] )
        , .SB_CORRECT(\SB_CORRECT[1][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C6 (.A_DOUT({nc2926, 
        nc2927, nc2928, nc2929, nc2930, nc2931, nc2932, nc2933, nc2934, 
        nc2935, nc2936, nc2937, nc2938, nc2939, nc2940, nc2941, nc2942, 
        nc2943, \R_DATA_TEMPR29[13] , \R_DATA_TEMPR29[12] }), .B_DOUT({
        nc2944, nc2945, nc2946, nc2947, nc2948, nc2949, nc2950, nc2951, 
        nc2952, nc2953, nc2954, nc2955, nc2956, nc2957, nc2958, nc2959, 
        nc2960, nc2961, nc2962, nc2963}), .DB_DETECT(
        \DB_DETECT[29][6] ), .SB_CORRECT(\SB_CORRECT[29][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0 (.A_DOUT({nc2964, 
        nc2965, nc2966, nc2967, nc2968, nc2969, nc2970, nc2971, nc2972, 
        nc2973, nc2974, nc2975, nc2976, nc2977, nc2978, nc2979, nc2980, 
        nc2981, \R_DATA_TEMPR23[1] , \R_DATA_TEMPR23[0] }), .B_DOUT({
        nc2982, nc2983, nc2984, nc2985, nc2986, nc2987, nc2988, nc2989, 
        nc2990, nc2991, nc2992, nc2993, nc2994, nc2995, nc2996, nc2997, 
        nc2998, nc2999, nc3000, nc3001}), .DB_DETECT(
        \DB_DETECT[23][0] ), .SB_CORRECT(\SB_CORRECT[23][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C10 (.A_DOUT({nc3002, 
        nc3003, nc3004, nc3005, nc3006, nc3007, nc3008, nc3009, nc3010, 
        nc3011, nc3012, nc3013, nc3014, nc3015, nc3016, nc3017, nc3018, 
        nc3019, \R_DATA_TEMPR0[21] , \R_DATA_TEMPR0[20] }), .B_DOUT({
        nc3020, nc3021, nc3022, nc3023, nc3024, nc3025, nc3026, nc3027, 
        nc3028, nc3029, nc3030, nc3031, nc3032, nc3033, nc3034, nc3035, 
        nc3036, nc3037, nc3038, nc3039}), .DB_DETECT(
        \DB_DETECT[0][10] ), .SB_CORRECT(\SB_CORRECT[0][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C4 (.A_DOUT({nc3040, 
        nc3041, nc3042, nc3043, nc3044, nc3045, nc3046, nc3047, nc3048, 
        nc3049, nc3050, nc3051, nc3052, nc3053, nc3054, nc3055, nc3056, 
        nc3057, \R_DATA_TEMPR18[9] , \R_DATA_TEMPR18[8] }), .B_DOUT({
        nc3058, nc3059, nc3060, nc3061, nc3062, nc3063, nc3064, nc3065, 
        nc3066, nc3067, nc3068, nc3069, nc3070, nc3071, nc3072, nc3073, 
        nc3074, nc3075, nc3076, nc3077}), .DB_DETECT(
        \DB_DETECT[18][4] ), .SB_CORRECT(\SB_CORRECT[18][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C7 (.A_DOUT({nc3078, 
        nc3079, nc3080, nc3081, nc3082, nc3083, nc3084, nc3085, nc3086, 
        nc3087, nc3088, nc3089, nc3090, nc3091, nc3092, nc3093, nc3094, 
        nc3095, \R_DATA_TEMPR20[15] , \R_DATA_TEMPR20[14] }), .B_DOUT({
        nc3096, nc3097, nc3098, nc3099, nc3100, nc3101, nc3102, nc3103, 
        nc3104, nc3105, nc3106, nc3107, nc3108, nc3109, nc3110, nc3111, 
        nc3112, nc3113, nc3114, nc3115}), .DB_DETECT(
        \DB_DETECT[20][7] ), .SB_CORRECT(\SB_CORRECT[20][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][7] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_232 (.A(\R_DATA_TEMPR0[20] ), .B(\R_DATA_TEMPR1[20] ), .C(
        \R_DATA_TEMPR2[20] ), .D(\R_DATA_TEMPR3[20] ), .Y(OR4_232_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C17 (.A_DOUT({
        nc3116, nc3117, nc3118, nc3119, nc3120, nc3121, nc3122, nc3123, 
        nc3124, nc3125, nc3126, nc3127, nc3128, nc3129, nc3130, nc3131, 
        nc3132, nc3133, \R_DATA_TEMPR28[35] , \R_DATA_TEMPR28[34] }), 
        .B_DOUT({nc3134, nc3135, nc3136, nc3137, nc3138, nc3139, 
        nc3140, nc3141, nc3142, nc3143, nc3144, nc3145, nc3146, nc3147, 
        nc3148, nc3149, nc3150, nc3151, nc3152, nc3153}), .DB_DETECT(
        \DB_DETECT[28][17] ), .SB_CORRECT(\SB_CORRECT[28][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[4]  (.A(CFG2_3_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[4] ));
    OR4 \OR4_R_DATA[15]  (.A(OR4_312_Y), .B(OR4_129_Y), .C(OR4_263_Y), 
        .D(OR4_156_Y), .Y(R_DATA[15]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C1 (.A_DOUT({nc3154, 
        nc3155, nc3156, nc3157, nc3158, nc3159, nc3160, nc3161, nc3162, 
        nc3163, nc3164, nc3165, nc3166, nc3167, nc3168, nc3169, nc3170, 
        nc3171, \R_DATA_TEMPR26[3] , \R_DATA_TEMPR26[2] }), .B_DOUT({
        nc3172, nc3173, nc3174, nc3175, nc3176, nc3177, nc3178, nc3179, 
        nc3180, nc3181, nc3182, nc3183, nc3184, nc3185, nc3186, nc3187, 
        nc3188, nc3189, nc3190, nc3191}), .DB_DETECT(
        \DB_DETECT[26][1] ), .SB_CORRECT(\SB_CORRECT[26][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C17 (.A_DOUT({nc3192, 
        nc3193, nc3194, nc3195, nc3196, nc3197, nc3198, nc3199, nc3200, 
        nc3201, nc3202, nc3203, nc3204, nc3205, nc3206, nc3207, nc3208, 
        nc3209, \R_DATA_TEMPR1[35] , \R_DATA_TEMPR1[34] }), .B_DOUT({
        nc3210, nc3211, nc3212, nc3213, nc3214, nc3215, nc3216, nc3217, 
        nc3218, nc3219, nc3220, nc3221, nc3222, nc3223, nc3224, nc3225, 
        nc3226, nc3227, nc3228, nc3229}), .DB_DETECT(
        \DB_DETECT[1][17] ), .SB_CORRECT(\SB_CORRECT[1][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_45 (.A(\R_DATA_TEMPR8[27] ), .B(\R_DATA_TEMPR9[27] ), .C(
        \R_DATA_TEMPR10[27] ), .D(\R_DATA_TEMPR11[27] ), .Y(OR4_45_Y));
    OR4 OR4_160 (.A(OR4_340_Y), .B(OR4_229_Y), .C(OR4_248_Y), .D(
        OR4_318_Y), .Y(OR4_160_Y));
    OR2 OR2_12 (.A(\R_DATA_TEMPR20[14] ), .B(\R_DATA_TEMPR21[14] ), .Y(
        OR2_12_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C6 (.A_DOUT({nc3230, 
        nc3231, nc3232, nc3233, nc3234, nc3235, nc3236, nc3237, nc3238, 
        nc3239, nc3240, nc3241, nc3242, nc3243, nc3244, nc3245, nc3246, 
        nc3247, \R_DATA_TEMPR15[13] , \R_DATA_TEMPR15[12] }), .B_DOUT({
        nc3248, nc3249, nc3250, nc3251, nc3252, nc3253, nc3254, nc3255, 
        nc3256, nc3257, nc3258, nc3259, nc3260, nc3261, nc3262, nc3263, 
        nc3264, nc3265, nc3266, nc3267}), .DB_DETECT(
        \DB_DETECT[15][6] ), .SB_CORRECT(\SB_CORRECT[15][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C5 (.A_DOUT({nc3268, 
        nc3269, nc3270, nc3271, nc3272, nc3273, nc3274, nc3275, nc3276, 
        nc3277, nc3278, nc3279, nc3280, nc3281, nc3282, nc3283, nc3284, 
        nc3285, \R_DATA_TEMPR22[11] , \R_DATA_TEMPR22[10] }), .B_DOUT({
        nc3286, nc3287, nc3288, nc3289, nc3290, nc3291, nc3292, nc3293, 
        nc3294, nc3295, nc3296, nc3297, nc3298, nc3299, nc3300, nc3301, 
        nc3302, nc3303, nc3304, nc3305}), .DB_DETECT(
        \DB_DETECT[22][5] ), .SB_CORRECT(\SB_CORRECT[22][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[23]  (.A(OR4_187_Y), .B(OR4_98_Y), .C(OR4_79_Y), 
        .D(OR4_68_Y), .Y(R_DATA[23]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C7 (.A_DOUT({nc3306, 
        nc3307, nc3308, nc3309, nc3310, nc3311, nc3312, nc3313, nc3314, 
        nc3315, nc3316, nc3317, nc3318, nc3319, nc3320, nc3321, nc3322, 
        nc3323, \R_DATA_TEMPR21[15] , \R_DATA_TEMPR21[14] }), .B_DOUT({
        nc3324, nc3325, nc3326, nc3327, nc3328, nc3329, nc3330, nc3331, 
        nc3332, nc3333, nc3334, nc3335, nc3336, nc3337, nc3338, nc3339, 
        nc3340, nc3341, nc3342, nc3343}), .DB_DETECT(
        \DB_DETECT[21][7] ), .SB_CORRECT(\SB_CORRECT[21][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][7] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_330 (.A(OR4_172_Y), .B(OR2_6_Y), .C(\R_DATA_TEMPR22[32] ), 
        .D(\R_DATA_TEMPR23[32] ), .Y(OR4_330_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C11 (.A_DOUT({nc3344, 
        nc3345, nc3346, nc3347, nc3348, nc3349, nc3350, nc3351, nc3352, 
        nc3353, nc3354, nc3355, nc3356, nc3357, nc3358, nc3359, nc3360, 
        nc3361, \R_DATA_TEMPR6[23] , \R_DATA_TEMPR6[22] }), .B_DOUT({
        nc3362, nc3363, nc3364, nc3365, nc3366, nc3367, nc3368, nc3369, 
        nc3370, nc3371, nc3372, nc3373, nc3374, nc3375, nc3376, nc3377, 
        nc3378, nc3379, nc3380, nc3381}), .DB_DETECT(
        \DB_DETECT[6][11] ), .SB_CORRECT(\SB_CORRECT[6][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1 (.A_DOUT({nc3382, 
        nc3383, nc3384, nc3385, nc3386, nc3387, nc3388, nc3389, nc3390, 
        nc3391, nc3392, nc3393, nc3394, nc3395, nc3396, nc3397, nc3398, 
        nc3399, \R_DATA_TEMPR10[3] , \R_DATA_TEMPR10[2] }), .B_DOUT({
        nc3400, nc3401, nc3402, nc3403, nc3404, nc3405, nc3406, nc3407, 
        nc3408, nc3409, nc3410, nc3411, nc3412, nc3413, nc3414, nc3415, 
        nc3416, nc3417, nc3418, nc3419}), .DB_DETECT(
        \DB_DETECT[10][1] ), .SB_CORRECT(\SB_CORRECT[10][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C8 (.A_DOUT({nc3420, 
        nc3421, nc3422, nc3423, nc3424, nc3425, nc3426, nc3427, nc3428, 
        nc3429, nc3430, nc3431, nc3432, nc3433, nc3434, nc3435, nc3436, 
        nc3437, \R_DATA_TEMPR28[17] , \R_DATA_TEMPR28[16] }), .B_DOUT({
        nc3438, nc3439, nc3440, nc3441, nc3442, nc3443, nc3444, nc3445, 
        nc3446, nc3447, nc3448, nc3449, nc3450, nc3451, nc3452, nc3453, 
        nc3454, nc3455, nc3456, nc3457}), .DB_DETECT(
        \DB_DETECT[28][8] ), .SB_CORRECT(\SB_CORRECT[28][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C12 (.A_DOUT({
        nc3458, nc3459, nc3460, nc3461, nc3462, nc3463, nc3464, nc3465, 
        nc3466, nc3467, nc3468, nc3469, nc3470, nc3471, nc3472, nc3473, 
        nc3474, nc3475, \R_DATA_TEMPR21[25] , \R_DATA_TEMPR21[24] }), 
        .B_DOUT({nc3476, nc3477, nc3478, nc3479, nc3480, nc3481, 
        nc3482, nc3483, nc3484, nc3485, nc3486, nc3487, nc3488, nc3489, 
        nc3490, nc3491, nc3492, nc3493, nc3494, nc3495}), .DB_DETECT(
        \DB_DETECT[21][12] ), .SB_CORRECT(\SB_CORRECT[21][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C18 (.A_DOUT({
        nc3496, nc3497, nc3498, nc3499, nc3500, nc3501, nc3502, nc3503, 
        nc3504, nc3505, nc3506, nc3507, nc3508, nc3509, nc3510, nc3511, 
        nc3512, nc3513, \R_DATA_TEMPR14[37] , \R_DATA_TEMPR14[36] }), 
        .B_DOUT({nc3514, nc3515, nc3516, nc3517, nc3518, nc3519, 
        nc3520, nc3521, nc3522, nc3523, nc3524, nc3525, nc3526, nc3527, 
        nc3528, nc3529, nc3530, nc3531, nc3532, nc3533}), .DB_DETECT(
        \DB_DETECT[14][18] ), .SB_CORRECT(\SB_CORRECT[14][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_287 (.A(\R_DATA_TEMPR0[0] ), .B(\R_DATA_TEMPR1[0] ), .C(
        \R_DATA_TEMPR2[0] ), .D(\R_DATA_TEMPR3[0] ), .Y(OR4_287_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C10 (.A_DOUT({
        nc3534, nc3535, nc3536, nc3537, nc3538, nc3539, nc3540, nc3541, 
        nc3542, nc3543, nc3544, nc3545, nc3546, nc3547, nc3548, nc3549, 
        nc3550, nc3551, \R_DATA_TEMPR21[21] , \R_DATA_TEMPR21[20] }), 
        .B_DOUT({nc3552, nc3553, nc3554, nc3555, nc3556, nc3557, 
        nc3558, nc3559, nc3560, nc3561, nc3562, nc3563, nc3564, nc3565, 
        nc3566, nc3567, nc3568, nc3569, nc3570, nc3571}), .DB_DETECT(
        \DB_DETECT[21][10] ), .SB_CORRECT(\SB_CORRECT[21][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_86 (.A(\R_DATA_TEMPR28[16] ), .B(\R_DATA_TEMPR29[16] ), .C(
        \R_DATA_TEMPR30[16] ), .D(\R_DATA_TEMPR31[16] ), .Y(OR4_86_Y));
    OR4 OR4_33 (.A(\R_DATA_TEMPR28[10] ), .B(\R_DATA_TEMPR29[10] ), .C(
        \R_DATA_TEMPR30[10] ), .D(\R_DATA_TEMPR31[10] ), .Y(OR4_33_Y));
    OR4 OR4_168 (.A(\R_DATA_TEMPR0[35] ), .B(\R_DATA_TEMPR1[35] ), .C(
        \R_DATA_TEMPR2[35] ), .D(\R_DATA_TEMPR3[35] ), .Y(OR4_168_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0 (.A_DOUT({nc3572, 
        nc3573, nc3574, nc3575, nc3576, nc3577, nc3578, nc3579, nc3580, 
        nc3581, nc3582, nc3583, nc3584, nc3585, nc3586, nc3587, nc3588, 
        nc3589, \R_DATA_TEMPR29[1] , \R_DATA_TEMPR29[0] }), .B_DOUT({
        nc3590, nc3591, nc3592, nc3593, nc3594, nc3595, nc3596, nc3597, 
        nc3598, nc3599, nc3600, nc3601, nc3602, nc3603, nc3604, nc3605, 
        nc3606, nc3607, nc3608, nc3609}), .DB_DETECT(
        \DB_DETECT[29][0] ), .SB_CORRECT(\SB_CORRECT[29][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1 (.A_DOUT({nc3610, 
        nc3611, nc3612, nc3613, nc3614, nc3615, nc3616, nc3617, nc3618, 
        nc3619, nc3620, nc3621, nc3622, nc3623, nc3624, nc3625, nc3626, 
        nc3627, \R_DATA_TEMPR8[3] , \R_DATA_TEMPR8[2] }), .B_DOUT({
        nc3628, nc3629, nc3630, nc3631, nc3632, nc3633, nc3634, nc3635, 
        nc3636, nc3637, nc3638, nc3639, nc3640, nc3641, nc3642, nc3643, 
        nc3644, nc3645, nc3646, nc3647}), .DB_DETECT(\DB_DETECT[8][1] )
        , .SB_CORRECT(\SB_CORRECT[8][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C14 (.A_DOUT({
        nc3648, nc3649, nc3650, nc3651, nc3652, nc3653, nc3654, nc3655, 
        nc3656, nc3657, nc3658, nc3659, nc3660, nc3661, nc3662, nc3663, 
        nc3664, nc3665, \R_DATA_TEMPR28[29] , \R_DATA_TEMPR28[28] }), 
        .B_DOUT({nc3666, nc3667, nc3668, nc3669, nc3670, nc3671, 
        nc3672, nc3673, nc3674, nc3675, nc3676, nc3677, nc3678, nc3679, 
        nc3680, nc3681, nc3682, nc3683, nc3684, nc3685}), .DB_DETECT(
        \DB_DETECT[28][14] ), .SB_CORRECT(\SB_CORRECT[28][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_187 (.A(OR4_305_Y), .B(OR4_233_Y), .C(OR4_227_Y), .D(
        OR4_93_Y), .Y(OR4_187_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C18 (.A_DOUT({
        nc3686, nc3687, nc3688, nc3689, nc3690, nc3691, nc3692, nc3693, 
        nc3694, nc3695, nc3696, nc3697, nc3698, nc3699, nc3700, nc3701, 
        nc3702, nc3703, \R_DATA_TEMPR15[37] , \R_DATA_TEMPR15[36] }), 
        .B_DOUT({nc3704, nc3705, nc3706, nc3707, nc3708, nc3709, 
        nc3710, nc3711, nc3712, nc3713, nc3714, nc3715, nc3716, nc3717, 
        nc3718, nc3719, nc3720, nc3721, nc3722, nc3723}), .DB_DETECT(
        \DB_DETECT[15][18] ), .SB_CORRECT(\SB_CORRECT[15][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_212 (.A(OR4_336_Y), .B(OR4_268_Y), .C(OR4_258_Y), .D(
        OR4_126_Y), .Y(OR4_212_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C16 (.A_DOUT({
        nc3724, nc3725, nc3726, nc3727, nc3728, nc3729, nc3730, nc3731, 
        nc3732, nc3733, nc3734, nc3735, nc3736, nc3737, nc3738, nc3739, 
        nc3740, nc3741, \R_DATA_TEMPR11[33] , \R_DATA_TEMPR11[32] }), 
        .B_DOUT({nc3742, nc3743, nc3744, nc3745, nc3746, nc3747, 
        nc3748, nc3749, nc3750, nc3751, nc3752, nc3753, nc3754, nc3755, 
        nc3756, nc3757, nc3758, nc3759, nc3760, nc3761}), .DB_DETECT(
        \DB_DETECT[11][16] ), .SB_CORRECT(\SB_CORRECT[11][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_353 (.A(\R_DATA_TEMPR12[0] ), .B(\R_DATA_TEMPR13[0] ), .C(
        \R_DATA_TEMPR14[0] ), .D(\R_DATA_TEMPR15[0] ), .Y(OR4_353_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C19 (.A_DOUT({
        nc3762, nc3763, nc3764, nc3765, nc3766, nc3767, nc3768, nc3769, 
        nc3770, nc3771, nc3772, nc3773, nc3774, nc3775, nc3776, nc3777, 
        nc3778, nc3779, \R_DATA_TEMPR17[39] , \R_DATA_TEMPR17[38] }), 
        .B_DOUT({nc3780, nc3781, nc3782, nc3783, nc3784, nc3785, 
        nc3786, nc3787, nc3788, nc3789, nc3790, nc3791, nc3792, nc3793, 
        nc3794, nc3795, nc3796, nc3797, nc3798, nc3799}), .DB_DETECT(
        \DB_DETECT[17][19] ), .SB_CORRECT(\SB_CORRECT[17][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C10 (.A_DOUT({
        nc3800, nc3801, nc3802, nc3803, nc3804, nc3805, nc3806, nc3807, 
        nc3808, nc3809, nc3810, nc3811, nc3812, nc3813, nc3814, nc3815, 
        nc3816, nc3817, \R_DATA_TEMPR13[21] , \R_DATA_TEMPR13[20] }), 
        .B_DOUT({nc3818, nc3819, nc3820, nc3821, nc3822, nc3823, 
        nc3824, nc3825, nc3826, nc3827, nc3828, nc3829, nc3830, nc3831, 
        nc3832, nc3833, nc3834, nc3835, nc3836, nc3837}), .DB_DETECT(
        \DB_DETECT[13][10] ), .SB_CORRECT(\SB_CORRECT[13][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C2 (.A_DOUT({nc3838, 
        nc3839, nc3840, nc3841, nc3842, nc3843, nc3844, nc3845, nc3846, 
        nc3847, nc3848, nc3849, nc3850, nc3851, nc3852, nc3853, nc3854, 
        nc3855, \R_DATA_TEMPR17[5] , \R_DATA_TEMPR17[4] }), .B_DOUT({
        nc3856, nc3857, nc3858, nc3859, nc3860, nc3861, nc3862, nc3863, 
        nc3864, nc3865, nc3866, nc3867, nc3868, nc3869, nc3870, nc3871, 
        nc3872, nc3873, nc3874, nc3875}), .DB_DETECT(
        \DB_DETECT[17][2] ), .SB_CORRECT(\SB_CORRECT[17][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C15 (.A_DOUT({
        nc3876, nc3877, nc3878, nc3879, nc3880, nc3881, nc3882, nc3883, 
        nc3884, nc3885, nc3886, nc3887, nc3888, nc3889, nc3890, nc3891, 
        nc3892, nc3893, \R_DATA_TEMPR13[31] , \R_DATA_TEMPR13[30] }), 
        .B_DOUT({nc3894, nc3895, nc3896, nc3897, nc3898, nc3899, 
        nc3900, nc3901, nc3902, nc3903, nc3904, nc3905, nc3906, nc3907, 
        nc3908, nc3909, nc3910, nc3911, nc3912, nc3913}), .DB_DETECT(
        \DB_DETECT[13][15] ), .SB_CORRECT(\SB_CORRECT[13][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_310 (.A(OR4_198_Y), .B(OR4_131_Y), .C(OR4_65_Y), .D(
        OR4_85_Y), .Y(OR4_310_Y));
    OR4 OR4_284 (.A(\R_DATA_TEMPR16[24] ), .B(\R_DATA_TEMPR17[24] ), 
        .C(\R_DATA_TEMPR18[24] ), .D(\R_DATA_TEMPR19[24] ), .Y(
        OR4_284_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C17 (.A_DOUT({nc3914, 
        nc3915, nc3916, nc3917, nc3918, nc3919, nc3920, nc3921, nc3922, 
        nc3923, nc3924, nc3925, nc3926, nc3927, nc3928, nc3929, nc3930, 
        nc3931, \R_DATA_TEMPR8[35] , \R_DATA_TEMPR8[34] }), .B_DOUT({
        nc3932, nc3933, nc3934, nc3935, nc3936, nc3937, nc3938, nc3939, 
        nc3940, nc3941, nc3942, nc3943, nc3944, nc3945, nc3946, nc3947, 
        nc3948, nc3949, nc3950, nc3951}), .DB_DETECT(
        \DB_DETECT[8][17] ), .SB_CORRECT(\SB_CORRECT[8][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_5 (.A(\R_DATA_TEMPR0[34] ), .B(\R_DATA_TEMPR1[34] ), .C(
        \R_DATA_TEMPR2[34] ), .D(\R_DATA_TEMPR3[34] ), .Y(OR4_5_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C2 (.A_DOUT({nc3952, 
        nc3953, nc3954, nc3955, nc3956, nc3957, nc3958, nc3959, nc3960, 
        nc3961, nc3962, nc3963, nc3964, nc3965, nc3966, nc3967, nc3968, 
        nc3969, \R_DATA_TEMPR8[5] , \R_DATA_TEMPR8[4] }), .B_DOUT({
        nc3970, nc3971, nc3972, nc3973, nc3974, nc3975, nc3976, nc3977, 
        nc3978, nc3979, nc3980, nc3981, nc3982, nc3983, nc3984, nc3985, 
        nc3986, nc3987, nc3988, nc3989}), .DB_DETECT(\DB_DETECT[8][2] )
        , .SB_CORRECT(\SB_CORRECT[8][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_307 (.A(\R_DATA_TEMPR0[26] ), .B(\R_DATA_TEMPR1[26] ), .C(
        \R_DATA_TEMPR2[26] ), .D(\R_DATA_TEMPR3[26] ), .Y(OR4_307_Y));
    OR4 OR4_100 (.A(\R_DATA_TEMPR16[12] ), .B(\R_DATA_TEMPR17[12] ), 
        .C(\R_DATA_TEMPR18[12] ), .D(\R_DATA_TEMPR19[12] ), .Y(
        OR4_100_Y));
    OR4 OR4_99 (.A(\R_DATA_TEMPR28[37] ), .B(\R_DATA_TEMPR29[37] ), .C(
        \R_DATA_TEMPR30[37] ), .D(\R_DATA_TEMPR31[37] ), .Y(OR4_99_Y));
    OR4 OR4_156 (.A(\R_DATA_TEMPR28[15] ), .B(\R_DATA_TEMPR29[15] ), 
        .C(\R_DATA_TEMPR30[15] ), .D(\R_DATA_TEMPR31[15] ), .Y(
        OR4_156_Y));
    OR2 OR2_36 (.A(\R_DATA_TEMPR20[27] ), .B(\R_DATA_TEMPR21[27] ), .Y(
        OR2_36_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1 (.A_DOUT({nc3990, 
        nc3991, nc3992, nc3993, nc3994, nc3995, nc3996, nc3997, nc3998, 
        nc3999, nc4000, nc4001, nc4002, nc4003, nc4004, nc4005, nc4006, 
        nc4007, \R_DATA_TEMPR14[3] , \R_DATA_TEMPR14[2] }), .B_DOUT({
        nc4008, nc4009, nc4010, nc4011, nc4012, nc4013, nc4014, nc4015, 
        nc4016, nc4017, nc4018, nc4019, nc4020, nc4021, nc4022, nc4023, 
        nc4024, nc4025, nc4026, nc4027}), .DB_DETECT(
        \DB_DETECT[14][1] ), .SB_CORRECT(\SB_CORRECT[14][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_24 (.A(\R_DATA_TEMPR20[17] ), .B(\R_DATA_TEMPR21[17] ), .Y(
        OR2_24_Y));
    OR4 OR4_68 (.A(\R_DATA_TEMPR28[23] ), .B(\R_DATA_TEMPR29[23] ), .C(
        \R_DATA_TEMPR30[23] ), .D(\R_DATA_TEMPR31[23] ), .Y(OR4_68_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C5 (.A_DOUT({nc4028, 
        nc4029, nc4030, nc4031, nc4032, nc4033, nc4034, nc4035, nc4036, 
        nc4037, nc4038, nc4039, nc4040, nc4041, nc4042, nc4043, nc4044, 
        nc4045, \R_DATA_TEMPR17[11] , \R_DATA_TEMPR17[10] }), .B_DOUT({
        nc4046, nc4047, nc4048, nc4049, nc4050, nc4051, nc4052, nc4053, 
        nc4054, nc4055, nc4056, nc4057, nc4058, nc4059, nc4060, nc4061, 
        nc4062, nc4063, nc4064, nc4065}), .DB_DETECT(
        \DB_DETECT[17][5] ), .SB_CORRECT(\SB_CORRECT[17][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C8 (.A_DOUT({nc4066, 
        nc4067, nc4068, nc4069, nc4070, nc4071, nc4072, nc4073, nc4074, 
        nc4075, nc4076, nc4077, nc4078, nc4079, nc4080, nc4081, nc4082, 
        nc4083, \R_DATA_TEMPR15[17] , \R_DATA_TEMPR15[16] }), .B_DOUT({
        nc4084, nc4085, nc4086, nc4087, nc4088, nc4089, nc4090, nc4091, 
        nc4092, nc4093, nc4094, nc4095, nc4096, nc4097, nc4098, nc4099, 
        nc4100, nc4101, nc4102, nc4103}), .DB_DETECT(
        \DB_DETECT[15][8] ), .SB_CORRECT(\SB_CORRECT[15][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_170 (.A(OR4_240_Y), .B(OR2_23_Y), .C(\R_DATA_TEMPR22[2] ), 
        .D(\R_DATA_TEMPR23[2] ), .Y(OR4_170_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C6 (.A_DOUT({nc4104, 
        nc4105, nc4106, nc4107, nc4108, nc4109, nc4110, nc4111, nc4112, 
        nc4113, nc4114, nc4115, nc4116, nc4117, nc4118, nc4119, nc4120, 
        nc4121, \R_DATA_TEMPR28[13] , \R_DATA_TEMPR28[12] }), .B_DOUT({
        nc4122, nc4123, nc4124, nc4125, nc4126, nc4127, nc4128, nc4129, 
        nc4130, nc4131, nc4132, nc4133, nc4134, nc4135, nc4136, nc4137, 
        nc4138, nc4139, nc4140, nc4141}), .DB_DETECT(
        \DB_DETECT[28][6] ), .SB_CORRECT(\SB_CORRECT[28][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C10 (.A_DOUT({
        nc4142, nc4143, nc4144, nc4145, nc4146, nc4147, nc4148, nc4149, 
        nc4150, nc4151, nc4152, nc4153, nc4154, nc4155, nc4156, nc4157, 
        nc4158, nc4159, \R_DATA_TEMPR30[21] , \R_DATA_TEMPR30[20] }), 
        .B_DOUT({nc4160, nc4161, nc4162, nc4163, nc4164, nc4165, 
        nc4166, nc4167, nc4168, nc4169, nc4170, nc4171, nc4172, nc4173, 
        nc4174, nc4175, nc4176, nc4177, nc4178, nc4179}), .DB_DETECT(
        \DB_DETECT[30][10] ), .SB_CORRECT(\SB_CORRECT[30][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_31 (.A(\R_DATA_TEMPR12[36] ), .B(\R_DATA_TEMPR13[36] ), .C(
        \R_DATA_TEMPR14[36] ), .D(\R_DATA_TEMPR15[36] ), .Y(OR4_31_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C5 (.A_DOUT({nc4180, 
        nc4181, nc4182, nc4183, nc4184, nc4185, nc4186, nc4187, nc4188, 
        nc4189, nc4190, nc4191, nc4192, nc4193, nc4194, nc4195, nc4196, 
        nc4197, \R_DATA_TEMPR15[11] , \R_DATA_TEMPR15[10] }), .B_DOUT({
        nc4198, nc4199, nc4200, nc4201, nc4202, nc4203, nc4204, nc4205, 
        nc4206, nc4207, nc4208, nc4209, nc4210, nc4211, nc4212, nc4213, 
        nc4214, nc4215, nc4216, nc4217}), .DB_DETECT(
        \DB_DETECT[15][5] ), .SB_CORRECT(\SB_CORRECT[15][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C16 (.A_DOUT({nc4218, 
        nc4219, nc4220, nc4221, nc4222, nc4223, nc4224, nc4225, nc4226, 
        nc4227, nc4228, nc4229, nc4230, nc4231, nc4232, nc4233, nc4234, 
        nc4235, \R_DATA_TEMPR9[33] , \R_DATA_TEMPR9[32] }), .B_DOUT({
        nc4236, nc4237, nc4238, nc4239, nc4240, nc4241, nc4242, nc4243, 
        nc4244, nc4245, nc4246, nc4247, nc4248, nc4249, nc4250, nc4251, 
        nc4252, nc4253, nc4254, nc4255}), .DB_DETECT(
        \DB_DETECT[9][16] ), .SB_CORRECT(\SB_CORRECT[9][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[31]  (.A(OR4_83_Y), .B(OR4_61_Y), .C(OR4_70_Y), .D(
        OR4_321_Y), .Y(R_DATA[31]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1 (.A_DOUT({nc4256, 
        nc4257, nc4258, nc4259, nc4260, nc4261, nc4262, nc4263, nc4264, 
        nc4265, nc4266, nc4267, nc4268, nc4269, nc4270, nc4271, nc4272, 
        nc4273, \R_DATA_TEMPR15[3] , \R_DATA_TEMPR15[2] }), .B_DOUT({
        nc4274, nc4275, nc4276, nc4277, nc4278, nc4279, nc4280, nc4281, 
        nc4282, nc4283, nc4284, nc4285, nc4286, nc4287, nc4288, nc4289, 
        nc4290, nc4291, nc4292, nc4293}), .DB_DETECT(
        \DB_DETECT[15][1] ), .SB_CORRECT(\SB_CORRECT[15][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_243 (.A(\R_DATA_TEMPR24[2] ), .B(\R_DATA_TEMPR25[2] ), .C(
        \R_DATA_TEMPR26[2] ), .D(\R_DATA_TEMPR27[2] ), .Y(OR4_243_Y));
    OR4 OR4_358 (.A(\R_DATA_TEMPR8[30] ), .B(\R_DATA_TEMPR9[30] ), .C(
        \R_DATA_TEMPR10[30] ), .D(\R_DATA_TEMPR11[30] ), .Y(OR4_358_Y));
    OR4 OR4_80 (.A(\R_DATA_TEMPR4[34] ), .B(\R_DATA_TEMPR5[34] ), .C(
        \R_DATA_TEMPR6[34] ), .D(\R_DATA_TEMPR7[34] ), .Y(OR4_80_Y));
    OR4 OR4_191 (.A(\R_DATA_TEMPR24[33] ), .B(\R_DATA_TEMPR25[33] ), 
        .C(\R_DATA_TEMPR26[33] ), .D(\R_DATA_TEMPR27[33] ), .Y(
        OR4_191_Y));
    OR4 OR4_108 (.A(\R_DATA_TEMPR16[18] ), .B(\R_DATA_TEMPR17[18] ), 
        .C(\R_DATA_TEMPR18[18] ), .D(\R_DATA_TEMPR19[18] ), .Y(
        OR4_108_Y));
    OR4 OR4_1 (.A(\R_DATA_TEMPR24[24] ), .B(\R_DATA_TEMPR25[24] ), .C(
        \R_DATA_TEMPR26[24] ), .D(\R_DATA_TEMPR27[24] ), .Y(OR4_1_Y));
    OR4 OR4_87 (.A(\R_DATA_TEMPR12[6] ), .B(\R_DATA_TEMPR13[6] ), .C(
        \R_DATA_TEMPR14[6] ), .D(\R_DATA_TEMPR15[6] ), .Y(OR4_87_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C13 (.A_DOUT({
        nc4294, nc4295, nc4296, nc4297, nc4298, nc4299, nc4300, nc4301, 
        nc4302, nc4303, nc4304, nc4305, nc4306, nc4307, nc4308, nc4309, 
        nc4310, nc4311, \R_DATA_TEMPR11[27] , \R_DATA_TEMPR11[26] }), 
        .B_DOUT({nc4312, nc4313, nc4314, nc4315, nc4316, nc4317, 
        nc4318, nc4319, nc4320, nc4321, nc4322, nc4323, nc4324, nc4325, 
        nc4326, nc4327, nc4328, nc4329, nc4330, nc4331}), .DB_DETECT(
        \DB_DETECT[11][13] ), .SB_CORRECT(\SB_CORRECT[11][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[30]  (.A(OR4_14_Y), .B(OR4_103_Y), .C(OR4_259_Y), 
        .D(OR4_128_Y), .Y(R_DATA[30]));
    OR4 OR4_178 (.A(\R_DATA_TEMPR4[11] ), .B(\R_DATA_TEMPR5[11] ), .C(
        \R_DATA_TEMPR6[11] ), .D(\R_DATA_TEMPR7[11] ), .Y(OR4_178_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C13 (.A_DOUT({nc4332, 
        nc4333, nc4334, nc4335, nc4336, nc4337, nc4338, nc4339, nc4340, 
        nc4341, nc4342, nc4343, nc4344, nc4345, nc4346, nc4347, nc4348, 
        nc4349, \R_DATA_TEMPR1[27] , \R_DATA_TEMPR1[26] }), .B_DOUT({
        nc4350, nc4351, nc4352, nc4353, nc4354, nc4355, nc4356, nc4357, 
        nc4358, nc4359, nc4360, nc4361, nc4362, nc4363, nc4364, nc4365, 
        nc4366, nc4367, nc4368, nc4369}), .DB_DETECT(
        \DB_DETECT[1][13] ), .SB_CORRECT(\SB_CORRECT[1][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C1 (.A_DOUT({nc4370, 
        nc4371, nc4372, nc4373, nc4374, nc4375, nc4376, nc4377, nc4378, 
        nc4379, nc4380, nc4381, nc4382, nc4383, nc4384, nc4385, nc4386, 
        nc4387, \R_DATA_TEMPR27[3] , \R_DATA_TEMPR27[2] }), .B_DOUT({
        nc4388, nc4389, nc4390, nc4391, nc4392, nc4393, nc4394, nc4395, 
        nc4396, nc4397, nc4398, nc4399, nc4400, nc4401, nc4402, nc4403, 
        nc4404, nc4405, nc4406, nc4407}), .DB_DETECT(
        \DB_DETECT[27][1] ), .SB_CORRECT(\SB_CORRECT[27][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0 (.A_DOUT({nc4408, 
        nc4409, nc4410, nc4411, nc4412, nc4413, nc4414, nc4415, nc4416, 
        nc4417, nc4418, nc4419, nc4420, nc4421, nc4422, nc4423, nc4424, 
        nc4425, \R_DATA_TEMPR20[1] , \R_DATA_TEMPR20[0] }), .B_DOUT({
        nc4426, nc4427, nc4428, nc4429, nc4430, nc4431, nc4432, nc4433, 
        nc4434, nc4435, nc4436, nc4437, nc4438, nc4439, nc4440, nc4441, 
        nc4442, nc4443, nc4444, nc4445}), .DB_DETECT(
        \DB_DETECT[20][0] ), .SB_CORRECT(\SB_CORRECT[20][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C6 (.A_DOUT({nc4446, 
        nc4447, nc4448, nc4449, nc4450, nc4451, nc4452, nc4453, nc4454, 
        nc4455, nc4456, nc4457, nc4458, nc4459, nc4460, nc4461, nc4462, 
        nc4463, \R_DATA_TEMPR16[13] , \R_DATA_TEMPR16[12] }), .B_DOUT({
        nc4464, nc4465, nc4466, nc4467, nc4468, nc4469, nc4470, nc4471, 
        nc4472, nc4473, nc4474, nc4475, nc4476, nc4477, nc4478, nc4479, 
        nc4480, nc4481, nc4482, nc4483}), .DB_DETECT(
        \DB_DETECT[16][6] ), .SB_CORRECT(\SB_CORRECT[16][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C19 (.A_DOUT({
        nc4484, nc4485, nc4486, nc4487, nc4488, nc4489, nc4490, nc4491, 
        nc4492, nc4493, nc4494, nc4495, nc4496, nc4497, nc4498, nc4499, 
        nc4500, nc4501, \R_DATA_TEMPR12[39] , \R_DATA_TEMPR12[38] }), 
        .B_DOUT({nc4502, nc4503, nc4504, nc4505, nc4506, nc4507, 
        nc4508, nc4509, nc4510, nc4511, nc4512, nc4513, nc4514, nc4515, 
        nc4516, nc4517, nc4518, nc4519, nc4520, nc4521}), .DB_DETECT(
        \DB_DETECT[12][19] ), .SB_CORRECT(\SB_CORRECT[12][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_159 (.A(\R_DATA_TEMPR8[37] ), .B(\R_DATA_TEMPR9[37] ), .C(
        \R_DATA_TEMPR10[37] ), .D(\R_DATA_TEMPR11[37] ), .Y(OR4_159_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C2 (.A_DOUT({nc4522, 
        nc4523, nc4524, nc4525, nc4526, nc4527, nc4528, nc4529, nc4530, 
        nc4531, nc4532, nc4533, nc4534, nc4535, nc4536, nc4537, nc4538, 
        nc4539, \R_DATA_TEMPR15[5] , \R_DATA_TEMPR15[4] }), .B_DOUT({
        nc4540, nc4541, nc4542, nc4543, nc4544, nc4545, nc4546, nc4547, 
        nc4548, nc4549, nc4550, nc4551, nc4552, nc4553, nc4554, nc4555, 
        nc4556, nc4557, nc4558, nc4559}), .DB_DETECT(
        \DB_DETECT[15][2] ), .SB_CORRECT(\SB_CORRECT[15][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_165 (.A(\R_DATA_TEMPR16[31] ), .B(\R_DATA_TEMPR17[31] ), 
        .C(\R_DATA_TEMPR18[31] ), .D(\R_DATA_TEMPR19[31] ), .Y(
        OR4_165_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C12 (.A_DOUT({nc4560, 
        nc4561, nc4562, nc4563, nc4564, nc4565, nc4566, nc4567, nc4568, 
        nc4569, nc4570, nc4571, nc4572, nc4573, nc4574, nc4575, nc4576, 
        nc4577, \R_DATA_TEMPR4[25] , \R_DATA_TEMPR4[24] }), .B_DOUT({
        nc4578, nc4579, nc4580, nc4581, nc4582, nc4583, nc4584, nc4585, 
        nc4586, nc4587, nc4588, nc4589, nc4590, nc4591, nc4592, nc4593, 
        nc4594, nc4595, nc4596, nc4597}), .DB_DETECT(
        \DB_DETECT[4][12] ), .SB_CORRECT(\SB_CORRECT[4][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_133 (.A(\R_DATA_TEMPR28[25] ), .B(\R_DATA_TEMPR29[25] ), 
        .C(\R_DATA_TEMPR30[25] ), .D(\R_DATA_TEMPR31[25] ), .Y(
        OR4_133_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C13 (.A_DOUT({
        nc4598, nc4599, nc4600, nc4601, nc4602, nc4603, nc4604, nc4605, 
        nc4606, nc4607, nc4608, nc4609, nc4610, nc4611, nc4612, nc4613, 
        nc4614, nc4615, \R_DATA_TEMPR28[27] , \R_DATA_TEMPR28[26] }), 
        .B_DOUT({nc4616, nc4617, nc4618, nc4619, nc4620, nc4621, 
        nc4622, nc4623, nc4624, nc4625, nc4626, nc4627, nc4628, nc4629, 
        nc4630, nc4631, nc4632, nc4633, nc4634, nc4635}), .DB_DETECT(
        \DB_DETECT[28][13] ), .SB_CORRECT(\SB_CORRECT[28][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_92 (.A(\R_DATA_TEMPR16[11] ), .B(\R_DATA_TEMPR17[11] ), .C(
        \R_DATA_TEMPR18[11] ), .D(\R_DATA_TEMPR19[11] ), .Y(OR4_92_Y));
    OR4 \OR4_R_DATA[36]  (.A(OR4_246_Y), .B(OR4_88_Y), .C(OR4_142_Y), 
        .D(OR4_162_Y), .Y(R_DATA[36]));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[1]  (.A(CFG2_6_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[1] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C9 (.A_DOUT({nc4636, 
        nc4637, nc4638, nc4639, nc4640, nc4641, nc4642, nc4643, nc4644, 
        nc4645, nc4646, nc4647, nc4648, nc4649, nc4650, nc4651, nc4652, 
        nc4653, \R_DATA_TEMPR27[19] , \R_DATA_TEMPR27[18] }), .B_DOUT({
        nc4654, nc4655, nc4656, nc4657, nc4658, nc4659, nc4660, nc4661, 
        nc4662, nc4663, nc4664, nc4665, nc4666, nc4667, nc4668, nc4669, 
        nc4670, nc4671, nc4672, nc4673}), .DB_DETECT(
        \DB_DETECT[27][9] ), .SB_CORRECT(\SB_CORRECT[27][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0 (.A_DOUT({nc4674, 
        nc4675, nc4676, nc4677, nc4678, nc4679, nc4680, nc4681, nc4682, 
        nc4683, nc4684, nc4685, nc4686, nc4687, nc4688, nc4689, nc4690, 
        nc4691, \R_DATA_TEMPR8[1] , \R_DATA_TEMPR8[0] }), .B_DOUT({
        nc4692, nc4693, nc4694, nc4695, nc4696, nc4697, nc4698, nc4699, 
        nc4700, nc4701, nc4702, nc4703, nc4704, nc4705, nc4706, nc4707, 
        nc4708, nc4709, nc4710, nc4711}), .DB_DETECT(\DB_DETECT[8][0] )
        , .SB_CORRECT(\SB_CORRECT[8][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C4 (.A_DOUT({nc4712, 
        nc4713, nc4714, nc4715, nc4716, nc4717, nc4718, nc4719, nc4720, 
        nc4721, nc4722, nc4723, nc4724, nc4725, nc4726, nc4727, nc4728, 
        nc4729, \R_DATA_TEMPR23[9] , \R_DATA_TEMPR23[8] }), .B_DOUT({
        nc4730, nc4731, nc4732, nc4733, nc4734, nc4735, nc4736, nc4737, 
        nc4738, nc4739, nc4740, nc4741, nc4742, nc4743, nc4744, nc4745, 
        nc4746, nc4747, nc4748, nc4749}), .DB_DETECT(
        \DB_DETECT[23][4] ), .SB_CORRECT(\SB_CORRECT[23][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C17 (.A_DOUT({
        nc4750, nc4751, nc4752, nc4753, nc4754, nc4755, nc4756, nc4757, 
        nc4758, nc4759, nc4760, nc4761, nc4762, nc4763, nc4764, nc4765, 
        nc4766, nc4767, \R_DATA_TEMPR21[35] , \R_DATA_TEMPR21[34] }), 
        .B_DOUT({nc4768, nc4769, nc4770, nc4771, nc4772, nc4773, 
        nc4774, nc4775, nc4776, nc4777, nc4778, nc4779, nc4780, nc4781, 
        nc4782, nc4783, nc4784, nc4785, nc4786, nc4787}), .DB_DETECT(
        \DB_DETECT[21][17] ), .SB_CORRECT(\SB_CORRECT[21][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C3 (.A_DOUT({nc4788, 
        nc4789, nc4790, nc4791, nc4792, nc4793, nc4794, nc4795, nc4796, 
        nc4797, nc4798, nc4799, nc4800, nc4801, nc4802, nc4803, nc4804, 
        nc4805, \R_DATA_TEMPR25[7] , \R_DATA_TEMPR25[6] }), .B_DOUT({
        nc4806, nc4807, nc4808, nc4809, nc4810, nc4811, nc4812, nc4813, 
        nc4814, nc4815, nc4816, nc4817, nc4818, nc4819, nc4820, nc4821, 
        nc4822, nc4823, nc4824, nc4825}), .DB_DETECT(
        \DB_DETECT[25][3] ), .SB_CORRECT(\SB_CORRECT[25][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_30 (.A(\R_DATA_TEMPR20[37] ), .B(\R_DATA_TEMPR21[37] ), .Y(
        OR2_30_Y));
    CFG2 #( .INIT(4'h8) )  CFG2_0 (.A(W_ADDR[16]), .B(W_ADDR[15]), .Y(
        CFG2_0_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C10 (.A_DOUT({
        nc4826, nc4827, nc4828, nc4829, nc4830, nc4831, nc4832, nc4833, 
        nc4834, nc4835, nc4836, nc4837, nc4838, nc4839, nc4840, nc4841, 
        nc4842, nc4843, \R_DATA_TEMPR10[21] , \R_DATA_TEMPR10[20] }), 
        .B_DOUT({nc4844, nc4845, nc4846, nc4847, nc4848, nc4849, 
        nc4850, nc4851, nc4852, nc4853, nc4854, nc4855, nc4856, nc4857, 
        nc4858, nc4859, nc4860, nc4861, nc4862, nc4863}), .DB_DETECT(
        \DB_DETECT[10][10] ), .SB_CORRECT(\SB_CORRECT[10][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C4 (.A_DOUT({nc4864, 
        nc4865, nc4866, nc4867, nc4868, nc4869, nc4870, nc4871, nc4872, 
        nc4873, nc4874, nc4875, nc4876, nc4877, nc4878, nc4879, nc4880, 
        nc4881, \R_DATA_TEMPR20[9] , \R_DATA_TEMPR20[8] }), .B_DOUT({
        nc4882, nc4883, nc4884, nc4885, nc4886, nc4887, nc4888, nc4889, 
        nc4890, nc4891, nc4892, nc4893, nc4894, nc4895, nc4896, nc4897, 
        nc4898, nc4899, nc4900, nc4901}), .DB_DETECT(
        \DB_DETECT[20][4] ), .SB_CORRECT(\SB_CORRECT[20][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_324 (.A(\R_DATA_TEMPR0[12] ), .B(\R_DATA_TEMPR1[12] ), .C(
        \R_DATA_TEMPR2[12] ), .D(\R_DATA_TEMPR3[12] ), .Y(OR4_324_Y));
    OR4 OR4_265 (.A(\R_DATA_TEMPR8[31] ), .B(\R_DATA_TEMPR9[31] ), .C(
        \R_DATA_TEMPR10[31] ), .D(\R_DATA_TEMPR11[31] ), .Y(OR4_265_Y));
    OR4 OR4_49 (.A(\R_DATA_TEMPR16[26] ), .B(\R_DATA_TEMPR17[26] ), .C(
        \R_DATA_TEMPR18[26] ), .D(\R_DATA_TEMPR19[26] ), .Y(OR4_49_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C15 (.A_DOUT({
        nc4902, nc4903, nc4904, nc4905, nc4906, nc4907, nc4908, nc4909, 
        nc4910, nc4911, nc4912, nc4913, nc4914, nc4915, nc4916, nc4917, 
        nc4918, nc4919, \R_DATA_TEMPR10[31] , \R_DATA_TEMPR10[30] }), 
        .B_DOUT({nc4920, nc4921, nc4922, nc4923, nc4924, nc4925, 
        nc4926, nc4927, nc4928, nc4929, nc4930, nc4931, nc4932, nc4933, 
        nc4934, nc4935, nc4936, nc4937, nc4938, nc4939}), .DB_DETECT(
        \DB_DETECT[10][15] ), .SB_CORRECT(\SB_CORRECT[10][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_14 (.A(\R_DATA_TEMPR20[35] ), .B(\R_DATA_TEMPR21[35] ), .Y(
        OR2_14_Y));
    OR2 OR2_37 (.A(\R_DATA_TEMPR20[36] ), .B(\R_DATA_TEMPR21[36] ), .Y(
        OR2_37_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C8 (.A_DOUT({nc4940, 
        nc4941, nc4942, nc4943, nc4944, nc4945, nc4946, nc4947, nc4948, 
        nc4949, nc4950, nc4951, nc4952, nc4953, nc4954, nc4955, nc4956, 
        nc4957, \R_DATA_TEMPR26[17] , \R_DATA_TEMPR26[16] }), .B_DOUT({
        nc4958, nc4959, nc4960, nc4961, nc4962, nc4963, nc4964, nc4965, 
        nc4966, nc4967, nc4968, nc4969, nc4970, nc4971, nc4972, nc4973, 
        nc4974, nc4975, nc4976, nc4977}), .DB_DETECT(
        \DB_DETECT[26][8] ), .SB_CORRECT(\SB_CORRECT[26][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_121 (.A(\R_DATA_TEMPR24[4] ), .B(\R_DATA_TEMPR25[4] ), .C(
        \R_DATA_TEMPR26[4] ), .D(\R_DATA_TEMPR27[4] ), .Y(OR4_121_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0 (.A_DOUT({nc4978, 
        nc4979, nc4980, nc4981, nc4982, nc4983, nc4984, nc4985, nc4986, 
        nc4987, nc4988, nc4989, nc4990, nc4991, nc4992, nc4993, nc4994, 
        nc4995, \R_DATA_TEMPR4[1] , \R_DATA_TEMPR4[0] }), .B_DOUT({
        nc4996, nc4997, nc4998, nc4999, nc5000, nc5001, nc5002, nc5003, 
        nc5004, nc5005, nc5006, nc5007, nc5008, nc5009, nc5010, nc5011, 
        nc5012, nc5013, nc5014, nc5015}), .DB_DETECT(\DB_DETECT[4][0] )
        , .SB_CORRECT(\SB_CORRECT[4][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C7 (.A_DOUT({nc5016, 
        nc5017, nc5018, nc5019, nc5020, nc5021, nc5022, nc5023, nc5024, 
        nc5025, nc5026, nc5027, nc5028, nc5029, nc5030, nc5031, nc5032, 
        nc5033, \R_DATA_TEMPR28[15] , \R_DATA_TEMPR28[14] }), .B_DOUT({
        nc5034, nc5035, nc5036, nc5037, nc5038, nc5039, nc5040, nc5041, 
        nc5042, nc5043, nc5044, nc5045, nc5046, nc5047, nc5048, nc5049, 
        nc5050, nc5051, nc5052, nc5053}), .DB_DETECT(
        \DB_DETECT[28][7] ), .SB_CORRECT(\SB_CORRECT[28][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][7] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[18]  (.A(OR4_344_Y), .B(OR4_295_Y), .C(OR4_132_Y), 
        .D(OR4_173_Y), .Y(R_DATA[18]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C11 (.A_DOUT({
        nc5054, nc5055, nc5056, nc5057, nc5058, nc5059, nc5060, nc5061, 
        nc5062, nc5063, nc5064, nc5065, nc5066, nc5067, nc5068, nc5069, 
        nc5070, nc5071, \R_DATA_TEMPR16[23] , \R_DATA_TEMPR16[22] }), 
        .B_DOUT({nc5072, nc5073, nc5074, nc5075, nc5076, nc5077, 
        nc5078, nc5079, nc5080, nc5081, nc5082, nc5083, nc5084, nc5085, 
        nc5086, nc5087, nc5088, nc5089, nc5090, nc5091}), .DB_DETECT(
        \DB_DETECT[16][11] ), .SB_CORRECT(\SB_CORRECT[16][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C5 (.A_DOUT({nc5092, 
        nc5093, nc5094, nc5095, nc5096, nc5097, nc5098, nc5099, nc5100, 
        nc5101, nc5102, nc5103, nc5104, nc5105, nc5106, nc5107, nc5108, 
        nc5109, \R_DATA_TEMPR23[11] , \R_DATA_TEMPR23[10] }), .B_DOUT({
        nc5110, nc5111, nc5112, nc5113, nc5114, nc5115, nc5116, nc5117, 
        nc5118, nc5119, nc5120, nc5121, nc5122, nc5123, nc5124, nc5125, 
        nc5126, nc5127, nc5128, nc5129}), .DB_DETECT(
        \DB_DETECT[23][5] ), .SB_CORRECT(\SB_CORRECT[23][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C13 (.A_DOUT({nc5130, 
        nc5131, nc5132, nc5133, nc5134, nc5135, nc5136, nc5137, nc5138, 
        nc5139, nc5140, nc5141, nc5142, nc5143, nc5144, nc5145, nc5146, 
        nc5147, \R_DATA_TEMPR8[27] , \R_DATA_TEMPR8[26] }), .B_DOUT({
        nc5148, nc5149, nc5150, nc5151, nc5152, nc5153, nc5154, nc5155, 
        nc5156, nc5157, nc5158, nc5159, nc5160, nc5161, nc5162, nc5163, 
        nc5164, nc5165, nc5166, nc5167}), .DB_DETECT(
        \DB_DETECT[8][13] ), .SB_CORRECT(\SB_CORRECT[8][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_113 (.A(\R_DATA_TEMPR4[2] ), .B(\R_DATA_TEMPR5[2] ), .C(
        \R_DATA_TEMPR6[2] ), .D(\R_DATA_TEMPR7[2] ), .Y(OR4_113_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C15 (.A_DOUT({nc5168, 
        nc5169, nc5170, nc5171, nc5172, nc5173, nc5174, nc5175, nc5176, 
        nc5177, nc5178, nc5179, nc5180, nc5181, nc5182, nc5183, nc5184, 
        nc5185, \R_DATA_TEMPR6[31] , \R_DATA_TEMPR6[30] }), .B_DOUT({
        nc5186, nc5187, nc5188, nc5189, nc5190, nc5191, nc5192, nc5193, 
        nc5194, nc5195, nc5196, nc5197, nc5198, nc5199, nc5200, nc5201, 
        nc5202, nc5203, nc5204, nc5205}), .DB_DETECT(
        \DB_DETECT[6][15] ), .SB_CORRECT(\SB_CORRECT[6][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_132 (.A(\R_DATA_TEMPR24[18] ), .B(\R_DATA_TEMPR25[18] ), 
        .C(\R_DATA_TEMPR26[18] ), .D(\R_DATA_TEMPR27[18] ), .Y(
        OR4_132_Y));
    OR4 OR4_7 (.A(\R_DATA_TEMPR28[22] ), .B(\R_DATA_TEMPR29[22] ), .C(
        \R_DATA_TEMPR30[22] ), .D(\R_DATA_TEMPR31[22] ), .Y(OR4_7_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C16 (.A_DOUT({
        nc5206, nc5207, nc5208, nc5209, nc5210, nc5211, nc5212, nc5213, 
        nc5214, nc5215, nc5216, nc5217, nc5218, nc5219, nc5220, nc5221, 
        nc5222, nc5223, \R_DATA_TEMPR28[33] , \R_DATA_TEMPR28[32] }), 
        .B_DOUT({nc5224, nc5225, nc5226, nc5227, nc5228, nc5229, 
        nc5230, nc5231, nc5232, nc5233, nc5234, nc5235, nc5236, nc5237, 
        nc5238, nc5239, nc5240, nc5241, nc5242, nc5243}), .DB_DETECT(
        \DB_DETECT[28][16] ), .SB_CORRECT(\SB_CORRECT[28][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0 (.A_DOUT({nc5244, 
        nc5245, nc5246, nc5247, nc5248, nc5249, nc5250, nc5251, nc5252, 
        nc5253, nc5254, nc5255, nc5256, nc5257, nc5258, nc5259, nc5260, 
        nc5261, \R_DATA_TEMPR16[1] , \R_DATA_TEMPR16[0] }), .B_DOUT({
        nc5262, nc5263, nc5264, nc5265, nc5266, nc5267, nc5268, nc5269, 
        nc5270, nc5271, nc5272, nc5273, nc5274, nc5275, nc5276, nc5277, 
        nc5278, nc5279, nc5280, nc5281}), .DB_DETECT(
        \DB_DETECT[16][0] ), .SB_CORRECT(\SB_CORRECT[16][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C1 (.A_DOUT({nc5282, 
        nc5283, nc5284, nc5285, nc5286, nc5287, nc5288, nc5289, nc5290, 
        nc5291, nc5292, nc5293, nc5294, nc5295, nc5296, nc5297, nc5298, 
        nc5299, \R_DATA_TEMPR22[3] , \R_DATA_TEMPR22[2] }), .B_DOUT({
        nc5300, nc5301, nc5302, nc5303, nc5304, nc5305, nc5306, nc5307, 
        nc5308, nc5309, nc5310, nc5311, nc5312, nc5313, nc5314, nc5315, 
        nc5316, nc5317, nc5318, nc5319}), .DB_DETECT(
        \DB_DETECT[22][1] ), .SB_CORRECT(\SB_CORRECT[22][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C14 (.A_DOUT({
        nc5320, nc5321, nc5322, nc5323, nc5324, nc5325, nc5326, nc5327, 
        nc5328, nc5329, nc5330, nc5331, nc5332, nc5333, nc5334, nc5335, 
        nc5336, nc5337, \R_DATA_TEMPR21[29] , \R_DATA_TEMPR21[28] }), 
        .B_DOUT({nc5338, nc5339, nc5340, nc5341, nc5342, nc5343, 
        nc5344, nc5345, nc5346, nc5347, nc5348, nc5349, nc5350, nc5351, 
        nc5352, nc5353, nc5354, nc5355, nc5356, nc5357}), .DB_DETECT(
        \DB_DETECT[21][14] ), .SB_CORRECT(\SB_CORRECT[21][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_268 (.A(\R_DATA_TEMPR4[13] ), .B(\R_DATA_TEMPR5[13] ), .C(
        \R_DATA_TEMPR6[13] ), .D(\R_DATA_TEMPR7[13] ), .Y(OR4_268_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C3 (.A_DOUT({nc5358, 
        nc5359, nc5360, nc5361, nc5362, nc5363, nc5364, nc5365, nc5366, 
        nc5367, nc5368, nc5369, nc5370, nc5371, nc5372, nc5373, nc5374, 
        nc5375, \R_DATA_TEMPR7[7] , \R_DATA_TEMPR7[6] }), .B_DOUT({
        nc5376, nc5377, nc5378, nc5379, nc5380, nc5381, nc5382, nc5383, 
        nc5384, nc5385, nc5386, nc5387, nc5388, nc5389, nc5390, nc5391, 
        nc5392, nc5393, nc5394, nc5395}), .DB_DETECT(\DB_DETECT[7][3] )
        , .SB_CORRECT(\SB_CORRECT[7][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_180 (.A(OR4_139_Y), .B(OR2_9_Y), .C(\R_DATA_TEMPR22[3] ), 
        .D(\R_DATA_TEMPR23[3] ), .Y(OR4_180_Y));
    OR4 OR4_105 (.A(\R_DATA_TEMPR24[28] ), .B(\R_DATA_TEMPR25[28] ), 
        .C(\R_DATA_TEMPR26[28] ), .D(\R_DATA_TEMPR27[28] ), .Y(
        OR4_105_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C15 (.A_DOUT({
        nc5396, nc5397, nc5398, nc5399, nc5400, nc5401, nc5402, nc5403, 
        nc5404, nc5405, nc5406, nc5407, nc5408, nc5409, nc5410, nc5411, 
        nc5412, nc5413, \R_DATA_TEMPR28[31] , \R_DATA_TEMPR28[30] }), 
        .B_DOUT({nc5414, nc5415, nc5416, nc5417, nc5418, nc5419, 
        nc5420, nc5421, nc5422, nc5423, nc5424, nc5425, nc5426, nc5427, 
        nc5428, nc5429, nc5430, nc5431, nc5432, nc5433}), .DB_DETECT(
        \DB_DETECT[28][15] ), .SB_CORRECT(\SB_CORRECT[28][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_175 (.A(\R_DATA_TEMPR8[38] ), .B(\R_DATA_TEMPR9[38] ), .C(
        \R_DATA_TEMPR10[38] ), .D(\R_DATA_TEMPR11[38] ), .Y(OR4_175_Y));
    OR4 OR4_239 (.A(\R_DATA_TEMPR4[38] ), .B(\R_DATA_TEMPR5[38] ), .C(
        \R_DATA_TEMPR6[38] ), .D(\R_DATA_TEMPR7[38] ), .Y(OR4_239_Y));
    OR4 OR4_42 (.A(\R_DATA_TEMPR0[32] ), .B(\R_DATA_TEMPR1[32] ), .C(
        \R_DATA_TEMPR2[32] ), .D(\R_DATA_TEMPR3[32] ), .Y(OR4_42_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C10 (.A_DOUT({
        nc5434, nc5435, nc5436, nc5437, nc5438, nc5439, nc5440, nc5441, 
        nc5442, nc5443, nc5444, nc5445, nc5446, nc5447, nc5448, nc5449, 
        nc5450, nc5451, \R_DATA_TEMPR14[21] , \R_DATA_TEMPR14[20] }), 
        .B_DOUT({nc5452, nc5453, nc5454, nc5455, nc5456, nc5457, 
        nc5458, nc5459, nc5460, nc5461, nc5462, nc5463, nc5464, nc5465, 
        nc5466, nc5467, nc5468, nc5469, nc5470, nc5471}), .DB_DETECT(
        \DB_DETECT[14][10] ), .SB_CORRECT(\SB_CORRECT[14][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C9 (.A_DOUT({nc5472, 
        nc5473, nc5474, nc5475, nc5476, nc5477, nc5478, nc5479, nc5480, 
        nc5481, nc5482, nc5483, nc5484, nc5485, nc5486, nc5487, nc5488, 
        nc5489, \R_DATA_TEMPR8[19] , \R_DATA_TEMPR8[18] }), .B_DOUT({
        nc5490, nc5491, nc5492, nc5493, nc5494, nc5495, nc5496, nc5497, 
        nc5498, nc5499, nc5500, nc5501, nc5502, nc5503, nc5504, nc5505, 
        nc5506, nc5507, nc5508, nc5509}), .DB_DETECT(\DB_DETECT[8][9] )
        , .SB_CORRECT(\SB_CORRECT[8][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C15 (.A_DOUT({
        nc5510, nc5511, nc5512, nc5513, nc5514, nc5515, nc5516, nc5517, 
        nc5518, nc5519, nc5520, nc5521, nc5522, nc5523, nc5524, nc5525, 
        nc5526, nc5527, \R_DATA_TEMPR14[31] , \R_DATA_TEMPR14[30] }), 
        .B_DOUT({nc5528, nc5529, nc5530, nc5531, nc5532, nc5533, 
        nc5534, nc5535, nc5536, nc5537, nc5538, nc5539, nc5540, nc5541, 
        nc5542, nc5543, nc5544, nc5545, nc5546, nc5547}), .DB_DETECT(
        \DB_DETECT[14][15] ), .SB_CORRECT(\SB_CORRECT[14][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C6 (.A_DOUT({nc5548, 
        nc5549, nc5550, nc5551, nc5552, nc5553, nc5554, nc5555, nc5556, 
        nc5557, nc5558, nc5559, nc5560, nc5561, nc5562, nc5563, nc5564, 
        nc5565, \R_DATA_TEMPR31[13] , \R_DATA_TEMPR31[12] }), .B_DOUT({
        nc5566, nc5567, nc5568, nc5569, nc5570, nc5571, nc5572, nc5573, 
        nc5574, nc5575, nc5576, nc5577, nc5578, nc5579, nc5580, nc5581, 
        nc5582, nc5583, nc5584, nc5585}), .DB_DETECT(
        \DB_DETECT[31][6] ), .SB_CORRECT(\SB_CORRECT[31][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0 (.A_DOUT({nc5586, 
        nc5587, nc5588, nc5589, nc5590, nc5591, nc5592, nc5593, nc5594, 
        nc5595, nc5596, nc5597, nc5598, nc5599, nc5600, nc5601, nc5602, 
        nc5603, \R_DATA_TEMPR9[1] , \R_DATA_TEMPR9[0] }), .B_DOUT({
        nc5604, nc5605, nc5606, nc5607, nc5608, nc5609, nc5610, nc5611, 
        nc5612, nc5613, nc5614, nc5615, nc5616, nc5617, nc5618, nc5619, 
        nc5620, nc5621, nc5622, nc5623}), .DB_DETECT(\DB_DETECT[9][0] )
        , .SB_CORRECT(\SB_CORRECT[9][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C7 (.A_DOUT({nc5624, 
        nc5625, nc5626, nc5627, nc5628, nc5629, nc5630, nc5631, nc5632, 
        nc5633, nc5634, nc5635, nc5636, nc5637, nc5638, nc5639, nc5640, 
        nc5641, \R_DATA_TEMPR25[15] , \R_DATA_TEMPR25[14] }), .B_DOUT({
        nc5642, nc5643, nc5644, nc5645, nc5646, nc5647, nc5648, nc5649, 
        nc5650, nc5651, nc5652, nc5653, nc5654, nc5655, nc5656, nc5657, 
        nc5658, nc5659, nc5660, nc5661}), .DB_DETECT(
        \DB_DETECT[25][7] ), .SB_CORRECT(\SB_CORRECT[25][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][7] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C7 (.A_DOUT({nc5662, 
        nc5663, nc5664, nc5665, nc5666, nc5667, nc5668, nc5669, nc5670, 
        nc5671, nc5672, nc5673, nc5674, nc5675, nc5676, nc5677, nc5678, 
        nc5679, \R_DATA_TEMPR14[15] , \R_DATA_TEMPR14[14] }), .B_DOUT({
        nc5680, nc5681, nc5682, nc5683, nc5684, nc5685, nc5686, nc5687, 
        nc5688, nc5689, nc5690, nc5691, nc5692, nc5693, nc5694, nc5695, 
        nc5696, nc5697, nc5698, nc5699}), .DB_DETECT(
        \DB_DETECT[14][7] ), .SB_CORRECT(\SB_CORRECT[14][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][7] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_88 (.A(OR4_164_Y), .B(OR2_37_Y), .C(\R_DATA_TEMPR22[36] ), 
        .D(\R_DATA_TEMPR23[36] ), .Y(OR4_88_Y));
    OR4 OR4_205 (.A(OR4_137_Y), .B(OR2_1_Y), .C(\R_DATA_TEMPR22[33] ), 
        .D(\R_DATA_TEMPR23[33] ), .Y(OR4_205_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C10 (.A_DOUT({
        nc5700, nc5701, nc5702, nc5703, nc5704, nc5705, nc5706, nc5707, 
        nc5708, nc5709, nc5710, nc5711, nc5712, nc5713, nc5714, nc5715, 
        nc5716, nc5717, \R_DATA_TEMPR15[21] , \R_DATA_TEMPR15[20] }), 
        .B_DOUT({nc5718, nc5719, nc5720, nc5721, nc5722, nc5723, 
        nc5724, nc5725, nc5726, nc5727, nc5728, nc5729, nc5730, nc5731, 
        nc5732, nc5733, nc5734, nc5735, nc5736, nc5737}), .DB_DETECT(
        \DB_DETECT[15][10] ), .SB_CORRECT(\SB_CORRECT[15][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_188 (.A(\R_DATA_TEMPR28[1] ), .B(\R_DATA_TEMPR29[1] ), .C(
        \R_DATA_TEMPR30[1] ), .D(\R_DATA_TEMPR31[1] ), .Y(OR4_188_Y));
    OR4 OR4_196 (.A(\R_DATA_TEMPR24[12] ), .B(\R_DATA_TEMPR25[12] ), 
        .C(\R_DATA_TEMPR26[12] ), .D(\R_DATA_TEMPR27[12] ), .Y(
        OR4_196_Y));
    OR4 OR4_112 (.A(\R_DATA_TEMPR12[5] ), .B(\R_DATA_TEMPR13[5] ), .C(
        \R_DATA_TEMPR14[5] ), .D(\R_DATA_TEMPR15[5] ), .Y(OR4_112_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C15 (.A_DOUT({
        nc5738, nc5739, nc5740, nc5741, nc5742, nc5743, nc5744, nc5745, 
        nc5746, nc5747, nc5748, nc5749, nc5750, nc5751, nc5752, nc5753, 
        nc5754, nc5755, \R_DATA_TEMPR15[31] , \R_DATA_TEMPR15[30] }), 
        .B_DOUT({nc5756, nc5757, nc5758, nc5759, nc5760, nc5761, 
        nc5762, nc5763, nc5764, nc5765, nc5766, nc5767, nc5768, nc5769, 
        nc5770, nc5771, nc5772, nc5773, nc5774, nc5775}), .DB_DETECT(
        \DB_DETECT[15][15] ), .SB_CORRECT(\SB_CORRECT[15][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0 (.A_DOUT({nc5776, 
        nc5777, nc5778, nc5779, nc5780, nc5781, nc5782, nc5783, nc5784, 
        nc5785, nc5786, nc5787, nc5788, nc5789, nc5790, nc5791, nc5792, 
        nc5793, \R_DATA_TEMPR2[1] , \R_DATA_TEMPR2[0] }), .B_DOUT({
        nc5794, nc5795, nc5796, nc5797, nc5798, nc5799, nc5800, nc5801, 
        nc5802, nc5803, nc5804, nc5805, nc5806, nc5807, nc5808, nc5809, 
        nc5810, nc5811, nc5812, nc5813}), .DB_DETECT(\DB_DETECT[2][0] )
        , .SB_CORRECT(\SB_CORRECT[2][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C5 (.A_DOUT({nc5814, 
        nc5815, nc5816, nc5817, nc5818, nc5819, nc5820, nc5821, nc5822, 
        nc5823, nc5824, nc5825, nc5826, nc5827, nc5828, nc5829, nc5830, 
        nc5831, \R_DATA_TEMPR3[11] , \R_DATA_TEMPR3[10] }), .B_DOUT({
        nc5832, nc5833, nc5834, nc5835, nc5836, nc5837, nc5838, nc5839, 
        nc5840, nc5841, nc5842, nc5843, nc5844, nc5845, nc5846, nc5847, 
        nc5848, nc5849, nc5850, nc5851}), .DB_DETECT(\DB_DETECT[3][5] )
        , .SB_CORRECT(\SB_CORRECT[3][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_275 (.A(\R_DATA_TEMPR4[25] ), .B(\R_DATA_TEMPR5[25] ), .C(
        \R_DATA_TEMPR6[25] ), .D(\R_DATA_TEMPR7[25] ), .Y(OR4_275_Y));
    OR4 \OR4_R_DATA[37]  (.A(OR4_153_Y), .B(OR4_329_Y), .C(OR4_56_Y), 
        .D(OR4_99_Y), .Y(R_DATA[37]));
    OR4 OR4_257 (.A(\R_DATA_TEMPR4[32] ), .B(\R_DATA_TEMPR5[32] ), .C(
        \R_DATA_TEMPR6[32] ), .D(\R_DATA_TEMPR7[32] ), .Y(OR4_257_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C3 (.A_DOUT({nc5852, 
        nc5853, nc5854, nc5855, nc5856, nc5857, nc5858, nc5859, nc5860, 
        nc5861, nc5862, nc5863, nc5864, nc5865, nc5866, nc5867, nc5868, 
        nc5869, \R_DATA_TEMPR26[7] , \R_DATA_TEMPR26[6] }), .B_DOUT({
        nc5870, nc5871, nc5872, nc5873, nc5874, nc5875, nc5876, nc5877, 
        nc5878, nc5879, nc5880, nc5881, nc5882, nc5883, nc5884, nc5885, 
        nc5886, nc5887, nc5888, nc5889}), .DB_DETECT(
        \DB_DETECT[26][3] ), .SB_CORRECT(\SB_CORRECT[26][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_157 (.A(\R_DATA_TEMPR0[5] ), .B(\R_DATA_TEMPR1[5] ), .C(
        \R_DATA_TEMPR2[5] ), .D(\R_DATA_TEMPR3[5] ), .Y(OR4_157_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C19 (.A_DOUT({nc5890, 
        nc5891, nc5892, nc5893, nc5894, nc5895, nc5896, nc5897, nc5898, 
        nc5899, nc5900, nc5901, nc5902, nc5903, nc5904, nc5905, nc5906, 
        nc5907, \R_DATA_TEMPR4[39] , \R_DATA_TEMPR4[38] }), .B_DOUT({
        nc5908, nc5909, nc5910, nc5911, nc5912, nc5913, nc5914, nc5915, 
        nc5916, nc5917, nc5918, nc5919, nc5920, nc5921, nc5922, nc5923, 
        nc5924, nc5925, nc5926, nc5927}), .DB_DETECT(
        \DB_DETECT[4][19] ), .SB_CORRECT(\SB_CORRECT[4][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_219 (.A(\R_DATA_TEMPR12[27] ), .B(\R_DATA_TEMPR13[27] ), 
        .C(\R_DATA_TEMPR14[27] ), .D(\R_DATA_TEMPR15[27] ), .Y(
        OR4_219_Y));
    OR4 OR4_208 (.A(\R_DATA_TEMPR24[38] ), .B(\R_DATA_TEMPR25[38] ), 
        .C(\R_DATA_TEMPR26[38] ), .D(\R_DATA_TEMPR27[38] ), .Y(
        OR4_208_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C9 (.A_DOUT({nc5928, 
        nc5929, nc5930, nc5931, nc5932, nc5933, nc5934, nc5935, nc5936, 
        nc5937, nc5938, nc5939, nc5940, nc5941, nc5942, nc5943, nc5944, 
        nc5945, \R_DATA_TEMPR19[19] , \R_DATA_TEMPR19[18] }), .B_DOUT({
        nc5946, nc5947, nc5948, nc5949, nc5950, nc5951, nc5952, nc5953, 
        nc5954, nc5955, nc5956, nc5957, nc5958, nc5959, nc5960, nc5961, 
        nc5962, nc5963, nc5964, nc5965}), .DB_DETECT(
        \DB_DETECT[19][9] ), .SB_CORRECT(\SB_CORRECT[19][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_323 (.A(\R_DATA_TEMPR12[31] ), .B(\R_DATA_TEMPR13[31] ), 
        .C(\R_DATA_TEMPR14[31] ), .D(\R_DATA_TEMPR15[31] ), .Y(
        OR4_323_Y));
    OR4 \OR4_R_DATA[19]  (.A(OR4_117_Y), .B(OR4_26_Y), .C(OR4_9_Y), .D(
        OR4_304_Y), .Y(R_DATA[19]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C3 (.A_DOUT({nc5966, 
        nc5967, nc5968, nc5969, nc5970, nc5971, nc5972, nc5973, nc5974, 
        nc5975, nc5976, nc5977, nc5978, nc5979, nc5980, nc5981, nc5982, 
        nc5983, \R_DATA_TEMPR20[7] , \R_DATA_TEMPR20[6] }), .B_DOUT({
        nc5984, nc5985, nc5986, nc5987, nc5988, nc5989, nc5990, nc5991, 
        nc5992, nc5993, nc5994, nc5995, nc5996, nc5997, nc5998, nc5999, 
        nc6000, nc6001, nc6002, nc6003}), .DB_DETECT(
        \DB_DETECT[20][3] ), .SB_CORRECT(\SB_CORRECT[20][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C3 (.A_DOUT({nc6004, 
        nc6005, nc6006, nc6007, nc6008, nc6009, nc6010, nc6011, nc6012, 
        nc6013, nc6014, nc6015, nc6016, nc6017, nc6018, nc6019, nc6020, 
        nc6021, \R_DATA_TEMPR23[7] , \R_DATA_TEMPR23[6] }), .B_DOUT({
        nc6022, nc6023, nc6024, nc6025, nc6026, nc6027, nc6028, nc6029, 
        nc6030, nc6031, nc6032, nc6033, nc6034, nc6035, nc6036, nc6037, 
        nc6038, nc6039, nc6040, nc6041}), .DB_DETECT(
        \DB_DETECT[23][3] ), .SB_CORRECT(\SB_CORRECT[23][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C14 (.A_DOUT({nc6042, 
        nc6043, nc6044, nc6045, nc6046, nc6047, nc6048, nc6049, nc6050, 
        nc6051, nc6052, nc6053, nc6054, nc6055, nc6056, nc6057, nc6058, 
        nc6059, \R_DATA_TEMPR9[29] , \R_DATA_TEMPR9[28] }), .B_DOUT({
        nc6060, nc6061, nc6062, nc6063, nc6064, nc6065, nc6066, nc6067, 
        nc6068, nc6069, nc6070, nc6071, nc6072, nc6073, nc6074, nc6075, 
        nc6076, nc6077, nc6078, nc6079}), .DB_DETECT(
        \DB_DETECT[9][14] ), .SB_CORRECT(\SB_CORRECT[9][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_38 (.A(\R_DATA_TEMPR20[13] ), .B(\R_DATA_TEMPR21[13] ), .Y(
        OR2_38_Y));
    OR4 OR4_278 (.A(OR4_35_Y), .B(OR4_111_Y), .C(OR4_39_Y), .D(
        OR4_226_Y), .Y(OR4_278_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C12 (.A_DOUT({nc6080, 
        nc6081, nc6082, nc6083, nc6084, nc6085, nc6086, nc6087, nc6088, 
        nc6089, nc6090, nc6091, nc6092, nc6093, nc6094, nc6095, nc6096, 
        nc6097, \R_DATA_TEMPR3[25] , \R_DATA_TEMPR3[24] }), .B_DOUT({
        nc6098, nc6099, nc6100, nc6101, nc6102, nc6103, nc6104, nc6105, 
        nc6106, nc6107, nc6108, nc6109, nc6110, nc6111, nc6112, nc6113, 
        nc6114, nc6115, nc6116, nc6117}), .DB_DETECT(
        \DB_DETECT[3][12] ), .SB_CORRECT(\SB_CORRECT[3][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C14 (.A_DOUT({
        nc6118, nc6119, nc6120, nc6121, nc6122, nc6123, nc6124, nc6125, 
        nc6126, nc6127, nc6128, nc6129, nc6130, nc6131, nc6132, nc6133, 
        nc6134, nc6135, \R_DATA_TEMPR30[29] , \R_DATA_TEMPR30[28] }), 
        .B_DOUT({nc6136, nc6137, nc6138, nc6139, nc6140, nc6141, 
        nc6142, nc6143, nc6144, nc6145, nc6146, nc6147, nc6148, nc6149, 
        nc6150, nc6151, nc6152, nc6153, nc6154, nc6155}), .DB_DETECT(
        \DB_DETECT[30][14] ), .SB_CORRECT(\SB_CORRECT[30][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C13 (.A_DOUT({
        nc6156, nc6157, nc6158, nc6159, nc6160, nc6161, nc6162, nc6163, 
        nc6164, nc6165, nc6166, nc6167, nc6168, nc6169, nc6170, nc6171, 
        nc6172, nc6173, \R_DATA_TEMPR21[27] , \R_DATA_TEMPR21[26] }), 
        .B_DOUT({nc6174, nc6175, nc6176, nc6177, nc6178, nc6179, 
        nc6180, nc6181, nc6182, nc6183, nc6184, nc6185, nc6186, nc6187, 
        nc6188, nc6189, nc6190, nc6191, nc6192, nc6193}), .DB_DETECT(
        \DB_DETECT[21][13] ), .SB_CORRECT(\SB_CORRECT[21][13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][13] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_199 (.A(\R_DATA_TEMPR4[26] ), .B(\R_DATA_TEMPR5[26] ), .C(
        \R_DATA_TEMPR6[26] ), .D(\R_DATA_TEMPR7[26] ), .Y(OR4_199_Y));
    OR4 OR4_23 (.A(\R_DATA_TEMPR24[14] ), .B(\R_DATA_TEMPR25[14] ), .C(
        \R_DATA_TEMPR26[14] ), .D(\R_DATA_TEMPR27[14] ), .Y(OR4_23_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C1 (.A_DOUT({nc6194, 
        nc6195, nc6196, nc6197, nc6198, nc6199, nc6200, nc6201, nc6202, 
        nc6203, nc6204, nc6205, nc6206, nc6207, nc6208, nc6209, nc6210, 
        nc6211, \R_DATA_TEMPR31[3] , \R_DATA_TEMPR31[2] }), .B_DOUT({
        nc6212, nc6213, nc6214, nc6215, nc6216, nc6217, nc6218, nc6219, 
        nc6220, nc6221, nc6222, nc6223, nc6224, nc6225, nc6226, nc6227, 
        nc6228, nc6229, nc6230, nc6231}), .DB_DETECT(
        \DB_DETECT[31][1] ), .SB_CORRECT(\SB_CORRECT[31][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_254 (.A(\R_DATA_TEMPR0[19] ), .B(\R_DATA_TEMPR1[19] ), .C(
        \R_DATA_TEMPR2[19] ), .D(\R_DATA_TEMPR3[19] ), .Y(OR4_254_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C2 (.A_DOUT({nc6232, 
        nc6233, nc6234, nc6235, nc6236, nc6237, nc6238, nc6239, nc6240, 
        nc6241, nc6242, nc6243, nc6244, nc6245, nc6246, nc6247, nc6248, 
        nc6249, \R_DATA_TEMPR21[5] , \R_DATA_TEMPR21[4] }), .B_DOUT({
        nc6250, nc6251, nc6252, nc6253, nc6254, nc6255, nc6256, nc6257, 
        nc6258, nc6259, nc6260, nc6261, nc6262, nc6263, nc6264, nc6265, 
        nc6266, nc6267, nc6268, nc6269}), .DB_DETECT(
        \DB_DETECT[21][2] ), .SB_CORRECT(\SB_CORRECT[21][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_262 (.A(OR4_232_Y), .B(OR4_154_Y), .C(OR4_238_Y), .D(
        OR4_37_Y), .Y(OR4_262_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C8 (.A_DOUT({nc6270, 
        nc6271, nc6272, nc6273, nc6274, nc6275, nc6276, nc6277, nc6278, 
        nc6279, nc6280, nc6281, nc6282, nc6283, nc6284, nc6285, nc6286, 
        nc6287, \R_DATA_TEMPR30[17] , \R_DATA_TEMPR30[16] }), .B_DOUT({
        nc6288, nc6289, nc6290, nc6291, nc6292, nc6293, nc6294, nc6295, 
        nc6296, nc6297, nc6298, nc6299, nc6300, nc6301, nc6302, nc6303, 
        nc6304, nc6305, nc6306, nc6307}), .DB_DETECT(
        \DB_DETECT[30][8] ), .SB_CORRECT(\SB_CORRECT[30][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C19 (.A_DOUT({
        nc6308, nc6309, nc6310, nc6311, nc6312, nc6313, nc6314, nc6315, 
        nc6316, nc6317, nc6318, nc6319, nc6320, nc6321, nc6322, nc6323, 
        nc6324, nc6325, \R_DATA_TEMPR19[39] , \R_DATA_TEMPR19[38] }), 
        .B_DOUT({nc6326, nc6327, nc6328, nc6329, nc6330, nc6331, 
        nc6332, nc6333, nc6334, nc6335, nc6336, nc6337, nc6338, nc6339, 
        nc6340, nc6341, nc6342, nc6343, nc6344, nc6345}), .DB_DETECT(
        \DB_DETECT[19][19] ), .SB_CORRECT(\SB_CORRECT[19][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_126 (.A(\R_DATA_TEMPR12[13] ), .B(\R_DATA_TEMPR13[13] ), 
        .C(\R_DATA_TEMPR14[13] ), .D(\R_DATA_TEMPR15[13] ), .Y(
        OR4_126_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C2 (.A_DOUT({nc6346, 
        nc6347, nc6348, nc6349, nc6350, nc6351, nc6352, nc6353, nc6354, 
        nc6355, nc6356, nc6357, nc6358, nc6359, nc6360, nc6361, nc6362, 
        nc6363, \R_DATA_TEMPR18[5] , \R_DATA_TEMPR18[4] }), .B_DOUT({
        nc6364, nc6365, nc6366, nc6367, nc6368, nc6369, nc6370, nc6371, 
        nc6372, nc6373, nc6374, nc6375, nc6376, nc6377, nc6378, nc6379, 
        nc6380, nc6381, nc6382, nc6383}), .DB_DETECT(
        \DB_DETECT[18][2] ), .SB_CORRECT(\SB_CORRECT[18][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_94 (.A(\R_DATA_TEMPR0[21] ), .B(\R_DATA_TEMPR1[21] ), .C(
        \R_DATA_TEMPR2[21] ), .D(\R_DATA_TEMPR3[21] ), .Y(OR4_94_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C11 (.A_DOUT({
        nc6384, nc6385, nc6386, nc6387, nc6388, nc6389, nc6390, nc6391, 
        nc6392, nc6393, nc6394, nc6395, nc6396, nc6397, nc6398, nc6399, 
        nc6400, nc6401, \R_DATA_TEMPR17[23] , \R_DATA_TEMPR17[22] }), 
        .B_DOUT({nc6402, nc6403, nc6404, nc6405, nc6406, nc6407, 
        nc6408, nc6409, nc6410, nc6411, nc6412, nc6413, nc6414, nc6415, 
        nc6416, nc6417, nc6418, nc6419, nc6420, nc6421}), .DB_DETECT(
        \DB_DETECT[17][11] ), .SB_CORRECT(\SB_CORRECT[17][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C10 (.A_DOUT({nc6422, 
        nc6423, nc6424, nc6425, nc6426, nc6427, nc6428, nc6429, nc6430, 
        nc6431, nc6432, nc6433, nc6434, nc6435, nc6436, nc6437, nc6438, 
        nc6439, \R_DATA_TEMPR6[21] , \R_DATA_TEMPR6[20] }), .B_DOUT({
        nc6440, nc6441, nc6442, nc6443, nc6444, nc6445, nc6446, nc6447, 
        nc6448, nc6449, nc6450, nc6451, nc6452, nc6453, nc6454, nc6455, 
        nc6456, nc6457, nc6458, nc6459}), .DB_DETECT(
        \DB_DETECT[6][10] ), .SB_CORRECT(\SB_CORRECT[6][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_65 (.A(\R_DATA_TEMPR8[28] ), .B(\R_DATA_TEMPR9[28] ), .C(
        \R_DATA_TEMPR10[28] ), .D(\R_DATA_TEMPR11[28] ), .Y(OR4_65_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C9 (.A_DOUT({nc6460, 
        nc6461, nc6462, nc6463, nc6464, nc6465, nc6466, nc6467, nc6468, 
        nc6469, nc6470, nc6471, nc6472, nc6473, nc6474, nc6475, nc6476, 
        nc6477, \R_DATA_TEMPR25[19] , \R_DATA_TEMPR25[18] }), .B_DOUT({
        nc6478, nc6479, nc6480, nc6481, nc6482, nc6483, nc6484, nc6485, 
        nc6486, nc6487, nc6488, nc6489, nc6490, nc6491, nc6492, nc6493, 
        nc6494, nc6495, nc6496, nc6497}), .DB_DETECT(
        \DB_DETECT[25][9] ), .SB_CORRECT(\SB_CORRECT[25][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_355 (.A(\R_DATA_TEMPR4[29] ), .B(\R_DATA_TEMPR5[29] ), .C(
        \R_DATA_TEMPR6[29] ), .D(\R_DATA_TEMPR7[29] ), .Y(OR4_355_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C16 (.A_DOUT({nc6498, 
        nc6499, nc6500, nc6501, nc6502, nc6503, nc6504, nc6505, nc6506, 
        nc6507, nc6508, nc6509, nc6510, nc6511, nc6512, nc6513, nc6514, 
        nc6515, \R_DATA_TEMPR2[33] , \R_DATA_TEMPR2[32] }), .B_DOUT({
        nc6516, nc6517, nc6518, nc6519, nc6520, nc6521, nc6522, nc6523, 
        nc6524, nc6525, nc6526, nc6527, nc6528, nc6529, nc6530, nc6531, 
        nc6532, nc6533, nc6534, nc6535}), .DB_DETECT(
        \DB_DETECT[2][16] ), .SB_CORRECT(\SB_CORRECT[2][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_344 (.A(OR4_228_Y), .B(OR4_150_Y), .C(OR4_102_Y), .D(
        OR4_120_Y), .Y(OR4_344_Y));
    OR4 OR4_328 (.A(OR4_94_Y), .B(OR4_146_Y), .C(OR4_145_Y), .D(
        OR4_207_Y), .Y(OR4_328_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C9 (.A_DOUT({nc6536, 
        nc6537, nc6538, nc6539, nc6540, nc6541, nc6542, nc6543, nc6544, 
        nc6545, nc6546, nc6547, nc6548, nc6549, nc6550, nc6551, nc6552, 
        nc6553, \R_DATA_TEMPR21[19] , \R_DATA_TEMPR21[18] }), .B_DOUT({
        nc6554, nc6555, nc6556, nc6557, nc6558, nc6559, nc6560, nc6561, 
        nc6562, nc6563, nc6564, nc6565, nc6566, nc6567, nc6568, nc6569, 
        nc6570, nc6571, nc6572, nc6573}), .DB_DETECT(
        \DB_DETECT[21][9] ), .SB_CORRECT(\SB_CORRECT[21][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_185 (.A(\R_DATA_TEMPR28[14] ), .B(\R_DATA_TEMPR29[14] ), 
        .C(\R_DATA_TEMPR30[14] ), .D(\R_DATA_TEMPR31[14] ), .Y(
        OR4_185_Y));
    OR4 OR4_141 (.A(\R_DATA_TEMPR24[20] ), .B(\R_DATA_TEMPR25[20] ), 
        .C(\R_DATA_TEMPR26[20] ), .D(\R_DATA_TEMPR27[20] ), .Y(
        OR4_141_Y));
    OR4 OR4_36 (.A(\R_DATA_TEMPR12[22] ), .B(\R_DATA_TEMPR13[22] ), .C(
        \R_DATA_TEMPR14[22] ), .D(\R_DATA_TEMPR15[22] ), .Y(OR4_36_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C9 (.A_DOUT({nc6574, 
        nc6575, nc6576, nc6577, nc6578, nc6579, nc6580, nc6581, nc6582, 
        nc6583, nc6584, nc6585, nc6586, nc6587, nc6588, nc6589, nc6590, 
        nc6591, \R_DATA_TEMPR18[19] , \R_DATA_TEMPR18[18] }), .B_DOUT({
        nc6592, nc6593, nc6594, nc6595, nc6596, nc6597, nc6598, nc6599, 
        nc6600, nc6601, nc6602, nc6603, nc6604, nc6605, nc6606, nc6607, 
        nc6608, nc6609, nc6610, nc6611}), .DB_DETECT(
        \DB_DETECT[18][9] ), .SB_CORRECT(\SB_CORRECT[18][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C12 (.A_DOUT({
        nc6612, nc6613, nc6614, nc6615, nc6616, nc6617, nc6618, nc6619, 
        nc6620, nc6621, nc6622, nc6623, nc6624, nc6625, nc6626, nc6627, 
        nc6628, nc6629, \R_DATA_TEMPR30[25] , \R_DATA_TEMPR30[24] }), 
        .B_DOUT({nc6630, nc6631, nc6632, nc6633, nc6634, nc6635, 
        nc6636, nc6637, nc6638, nc6639, nc6640, nc6641, nc6642, nc6643, 
        nc6644, nc6645, nc6646, nc6647, nc6648, nc6649}), .DB_DETECT(
        \DB_DETECT[30][12] ), .SB_CORRECT(\SB_CORRECT[30][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C18 (.A_DOUT({
        nc6650, nc6651, nc6652, nc6653, nc6654, nc6655, nc6656, nc6657, 
        nc6658, nc6659, nc6660, nc6661, nc6662, nc6663, nc6664, nc6665, 
        nc6666, nc6667, \R_DATA_TEMPR18[37] , \R_DATA_TEMPR18[36] }), 
        .B_DOUT({nc6668, nc6669, nc6670, nc6671, nc6672, nc6673, 
        nc6674, nc6675, nc6676, nc6677, nc6678, nc6679, nc6680, nc6681, 
        nc6682, nc6683, nc6684, nc6685, nc6686, nc6687}), .DB_DETECT(
        \DB_DETECT[18][18] ), .SB_CORRECT(\SB_CORRECT[18][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_21 (.A(\R_DATA_TEMPR16[23] ), .B(\R_DATA_TEMPR17[23] ), .C(
        \R_DATA_TEMPR18[23] ), .D(\R_DATA_TEMPR19[23] ), .Y(OR4_21_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C3 (.A_DOUT({nc6688, 
        nc6689, nc6690, nc6691, nc6692, nc6693, nc6694, nc6695, nc6696, 
        nc6697, nc6698, nc6699, nc6700, nc6701, nc6702, nc6703, nc6704, 
        nc6705, \R_DATA_TEMPR29[7] , \R_DATA_TEMPR29[6] }), .B_DOUT({
        nc6706, nc6707, nc6708, nc6709, nc6710, nc6711, nc6712, nc6713, 
        nc6714, nc6715, nc6716, nc6717, nc6718, nc6719, nc6720, nc6721, 
        nc6722, nc6723, nc6724, nc6725}), .DB_DETECT(
        \DB_DETECT[29][3] ), .SB_CORRECT(\SB_CORRECT[29][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C16 (.A_DOUT({
        nc6726, nc6727, nc6728, nc6729, nc6730, nc6731, nc6732, nc6733, 
        nc6734, nc6735, nc6736, nc6737, nc6738, nc6739, nc6740, nc6741, 
        nc6742, nc6743, \R_DATA_TEMPR21[33] , \R_DATA_TEMPR21[32] }), 
        .B_DOUT({nc6744, nc6745, nc6746, nc6747, nc6748, nc6749, 
        nc6750, nc6751, nc6752, nc6753, nc6754, nc6755, nc6756, nc6757, 
        nc6758, nc6759, nc6760, nc6761, nc6762, nc6763}), .DB_DETECT(
        \DB_DETECT[21][16] ), .SB_CORRECT(\SB_CORRECT[21][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[3]  (.A(CFG2_5_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[3] ));
    OR4 OR4_129 (.A(OR4_349_Y), .B(OR2_7_Y), .C(\R_DATA_TEMPR22[15] ), 
        .D(\R_DATA_TEMPR23[15] ), .Y(OR4_129_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C16 (.A_DOUT({nc6764, 
        nc6765, nc6766, nc6767, nc6768, nc6769, nc6770, nc6771, nc6772, 
        nc6773, nc6774, nc6775, nc6776, nc6777, nc6778, nc6779, nc6780, 
        nc6781, \R_DATA_TEMPR7[33] , \R_DATA_TEMPR7[32] }), .B_DOUT({
        nc6782, nc6783, nc6784, nc6785, nc6786, nc6787, nc6788, nc6789, 
        nc6790, nc6791, nc6792, nc6793, nc6794, nc6795, nc6796, nc6797, 
        nc6798, nc6799, nc6800, nc6801}), .DB_DETECT(
        \DB_DETECT[7][16] ), .SB_CORRECT(\SB_CORRECT[7][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0 (.A_DOUT({nc6802, 
        nc6803, nc6804, nc6805, nc6806, nc6807, nc6808, nc6809, nc6810, 
        nc6811, nc6812, nc6813, nc6814, nc6815, nc6816, nc6817, nc6818, 
        nc6819, \R_DATA_TEMPR24[1] , \R_DATA_TEMPR24[0] }), .B_DOUT({
        nc6820, nc6821, nc6822, nc6823, nc6824, nc6825, nc6826, nc6827, 
        nc6828, nc6829, nc6830, nc6831, nc6832, nc6833, nc6834, nc6835, 
        nc6836, nc6837, nc6838, nc6839}), .DB_DETECT(
        \DB_DETECT[24][0] ), .SB_CORRECT(\SB_CORRECT[24][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_285 (.A(OR4_59_Y), .B(OR4_275_Y), .C(OR4_290_Y), .D(
        OR4_115_Y), .Y(OR4_285_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C1 (.A_DOUT({nc6840, 
        nc6841, nc6842, nc6843, nc6844, nc6845, nc6846, nc6847, nc6848, 
        nc6849, nc6850, nc6851, nc6852, nc6853, nc6854, nc6855, nc6856, 
        nc6857, \R_DATA_TEMPR29[3] , \R_DATA_TEMPR29[2] }), .B_DOUT({
        nc6858, nc6859, nc6860, nc6861, nc6862, nc6863, nc6864, nc6865, 
        nc6866, nc6867, nc6868, nc6869, nc6870, nc6871, nc6872, nc6873, 
        nc6874, nc6875, nc6876, nc6877}), .DB_DETECT(
        \DB_DETECT[29][1] ), .SB_CORRECT(\SB_CORRECT[29][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C15 (.A_DOUT({
        nc6878, nc6879, nc6880, nc6881, nc6882, nc6883, nc6884, nc6885, 
        nc6886, nc6887, nc6888, nc6889, nc6890, nc6891, nc6892, nc6893, 
        nc6894, nc6895, \R_DATA_TEMPR21[31] , \R_DATA_TEMPR21[30] }), 
        .B_DOUT({nc6896, nc6897, nc6898, nc6899, nc6900, nc6901, 
        nc6902, nc6903, nc6904, nc6905, nc6906, nc6907, nc6908, nc6909, 
        nc6910, nc6911, nc6912, nc6913, nc6914, nc6915}), .DB_DETECT(
        \DB_DETECT[21][15] ), .SB_CORRECT(\SB_CORRECT[21][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C9 (.A_DOUT({nc6916, 
        nc6917, nc6918, nc6919, nc6920, nc6921, nc6922, nc6923, nc6924, 
        nc6925, nc6926, nc6927, nc6928, nc6929, nc6930, nc6931, nc6932, 
        nc6933, \R_DATA_TEMPR12[19] , \R_DATA_TEMPR12[18] }), .B_DOUT({
        nc6934, nc6935, nc6936, nc6937, nc6938, nc6939, nc6940, nc6941, 
        nc6942, nc6943, nc6944, nc6945, nc6946, nc6947, nc6948, nc6949, 
        nc6950, nc6951, nc6952, nc6953}), .DB_DETECT(
        \DB_DETECT[12][9] ), .SB_CORRECT(\SB_CORRECT[12][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_202 (.A(\R_DATA_TEMPR28[21] ), .B(\R_DATA_TEMPR29[21] ), 
        .C(\R_DATA_TEMPR30[21] ), .D(\R_DATA_TEMPR31[21] ), .Y(
        OR4_202_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C11 (.A_DOUT({
        nc6954, nc6955, nc6956, nc6957, nc6958, nc6959, nc6960, nc6961, 
        nc6962, nc6963, nc6964, nc6965, nc6966, nc6967, nc6968, nc6969, 
        nc6970, nc6971, \R_DATA_TEMPR12[23] , \R_DATA_TEMPR12[22] }), 
        .B_DOUT({nc6972, nc6973, nc6974, nc6975, nc6976, nc6977, 
        nc6978, nc6979, nc6980, nc6981, nc6982, nc6983, nc6984, nc6985, 
        nc6986, nc6987, nc6988, nc6989, nc6990, nc6991}), .DB_DETECT(
        \DB_DETECT[12][11] ), .SB_CORRECT(\SB_CORRECT[12][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_272 (.A(\R_DATA_TEMPR4[30] ), .B(\R_DATA_TEMPR5[30] ), .C(
        \R_DATA_TEMPR6[30] ), .D(\R_DATA_TEMPR7[30] ), .Y(OR4_272_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C18 (.A_DOUT({nc6992, 
        nc6993, nc6994, nc6995, nc6996, nc6997, nc6998, nc6999, nc7000, 
        nc7001, nc7002, nc7003, nc7004, nc7005, nc7006, nc7007, nc7008, 
        nc7009, \R_DATA_TEMPR9[37] , \R_DATA_TEMPR9[36] }), .B_DOUT({
        nc7010, nc7011, nc7012, nc7013, nc7014, nc7015, nc7016, nc7017, 
        nc7018, nc7019, nc7020, nc7021, nc7022, nc7023, nc7024, nc7025, 
        nc7026, nc7027, nc7028, nc7029}), .DB_DETECT(
        \DB_DETECT[9][18] ), .SB_CORRECT(\SB_CORRECT[9][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C8 (.A_DOUT({nc7030, 
        nc7031, nc7032, nc7033, nc7034, nc7035, nc7036, nc7037, nc7038, 
        nc7039, nc7040, nc7041, nc7042, nc7043, nc7044, nc7045, nc7046, 
        nc7047, \R_DATA_TEMPR21[17] , \R_DATA_TEMPR21[16] }), .B_DOUT({
        nc7048, nc7049, nc7050, nc7051, nc7052, nc7053, nc7054, nc7055, 
        nc7056, nc7057, nc7058, nc7059, nc7060, nc7061, nc7062, nc7063, 
        nc7064, nc7065, nc7066, nc7067}), .DB_DETECT(
        \DB_DETECT[21][8] ), .SB_CORRECT(\SB_CORRECT[21][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_44 (.A(\R_DATA_TEMPR4[7] ), .B(\R_DATA_TEMPR5[7] ), .C(
        \R_DATA_TEMPR6[7] ), .D(\R_DATA_TEMPR7[7] ), .Y(OR4_44_Y));
    OR4 OR4_300 (.A(\R_DATA_TEMPR12[14] ), .B(\R_DATA_TEMPR13[14] ), 
        .C(\R_DATA_TEMPR14[14] ), .D(\R_DATA_TEMPR15[14] ), .Y(
        OR4_300_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[0]  (.A(CFG2_4_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[0] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C8 (.A_DOUT({nc7068, 
        nc7069, nc7070, nc7071, nc7072, nc7073, nc7074, nc7075, nc7076, 
        nc7077, nc7078, nc7079, nc7080, nc7081, nc7082, nc7083, nc7084, 
        nc7085, \R_DATA_TEMPR14[17] , \R_DATA_TEMPR14[16] }), .B_DOUT({
        nc7086, nc7087, nc7088, nc7089, nc7090, nc7091, nc7092, nc7093, 
        nc7094, nc7095, nc7096, nc7097, nc7098, nc7099, nc7100, nc7101, 
        nc7102, nc7103, nc7104, nc7105}), .DB_DETECT(
        \DB_DETECT[14][8] ), .SB_CORRECT(\SB_CORRECT[14][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C14 (.A_DOUT({
        nc7106, nc7107, nc7108, nc7109, nc7110, nc7111, nc7112, nc7113, 
        nc7114, nc7115, nc7116, nc7117, nc7118, nc7119, nc7120, nc7121, 
        nc7122, nc7123, \R_DATA_TEMPR16[29] , \R_DATA_TEMPR16[28] }), 
        .B_DOUT({nc7124, nc7125, nc7126, nc7127, nc7128, nc7129, 
        nc7130, nc7131, nc7132, nc7133, nc7134, nc7135, nc7136, nc7137, 
        nc7138, nc7139, nc7140, nc7141, nc7142, nc7143}), .DB_DETECT(
        \DB_DETECT[16][14] ), .SB_CORRECT(\SB_CORRECT[16][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C4 (.A_DOUT({nc7144, 
        nc7145, nc7146, nc7147, nc7148, nc7149, nc7150, nc7151, nc7152, 
        nc7153, nc7154, nc7155, nc7156, nc7157, nc7158, nc7159, nc7160, 
        nc7161, \R_DATA_TEMPR17[9] , \R_DATA_TEMPR17[8] }), .B_DOUT({
        nc7162, nc7163, nc7164, nc7165, nc7166, nc7167, nc7168, nc7169, 
        nc7170, nc7171, nc7172, nc7173, nc7174, nc7175, nc7176, nc7177, 
        nc7178, nc7179, nc7180, nc7181}), .DB_DETECT(
        \DB_DETECT[17][4] ), .SB_CORRECT(\SB_CORRECT[17][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0 (.A_DOUT({nc7182, 
        nc7183, nc7184, nc7185, nc7186, nc7187, nc7188, nc7189, nc7190, 
        nc7191, nc7192, nc7193, nc7194, nc7195, nc7196, nc7197, nc7198, 
        nc7199, \R_DATA_TEMPR18[1] , \R_DATA_TEMPR18[0] }), .B_DOUT({
        nc7200, nc7201, nc7202, nc7203, nc7204, nc7205, nc7206, nc7207, 
        nc7208, nc7209, nc7210, nc7211, nc7212, nc7213, nc7214, nc7215, 
        nc7216, nc7217, nc7218, nc7219}), .DB_DETECT(
        \DB_DETECT[18][0] ), .SB_CORRECT(\SB_CORRECT[18][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C1 (.A_DOUT({nc7220, 
        nc7221, nc7222, nc7223, nc7224, nc7225, nc7226, nc7227, nc7228, 
        nc7229, nc7230, nc7231, nc7232, nc7233, nc7234, nc7235, nc7236, 
        nc7237, \R_DATA_TEMPR18[3] , \R_DATA_TEMPR18[2] }), .B_DOUT({
        nc7238, nc7239, nc7240, nc7241, nc7242, nc7243, nc7244, nc7245, 
        nc7246, nc7247, nc7248, nc7249, nc7250, nc7251, nc7252, nc7253, 
        nc7254, nc7255, nc7256, nc7257}), .DB_DETECT(
        \DB_DETECT[18][1] ), .SB_CORRECT(\SB_CORRECT[18][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_288 (.A(\R_DATA_TEMPR4[5] ), .B(\R_DATA_TEMPR5[5] ), .C(
        \R_DATA_TEMPR6[5] ), .D(\R_DATA_TEMPR7[5] ), .Y(OR4_288_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C2 (.A_DOUT({nc7258, 
        nc7259, nc7260, nc7261, nc7262, nc7263, nc7264, nc7265, nc7266, 
        nc7267, nc7268, nc7269, nc7270, nc7271, nc7272, nc7273, nc7274, 
        nc7275, \R_DATA_TEMPR29[5] , \R_DATA_TEMPR29[4] }), .B_DOUT({
        nc7276, nc7277, nc7278, nc7279, nc7280, nc7281, nc7282, nc7283, 
        nc7284, nc7285, nc7286, nc7287, nc7288, nc7289, nc7290, nc7291, 
        nc7292, nc7293, nc7294, nc7295}), .DB_DETECT(
        \DB_DETECT[29][2] ), .SB_CORRECT(\SB_CORRECT[29][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C16 (.A_DOUT({nc7296, 
        nc7297, nc7298, nc7299, nc7300, nc7301, nc7302, nc7303, nc7304, 
        nc7305, nc7306, nc7307, nc7308, nc7309, nc7310, nc7311, nc7312, 
        nc7313, \R_DATA_TEMPR5[33] , \R_DATA_TEMPR5[32] }), .B_DOUT({
        nc7314, nc7315, nc7316, nc7317, nc7318, nc7319, nc7320, nc7321, 
        nc7322, nc7323, nc7324, nc7325, nc7326, nc7327, nc7328, nc7329, 
        nc7330, nc7331, nc7332, nc7333}), .DB_DETECT(
        \DB_DETECT[5][16] ), .SB_CORRECT(\SB_CORRECT[5][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C17 (.A_DOUT({
        nc7334, nc7335, nc7336, nc7337, nc7338, nc7339, nc7340, nc7341, 
        nc7342, nc7343, nc7344, nc7345, nc7346, nc7347, nc7348, nc7349, 
        nc7350, nc7351, \R_DATA_TEMPR13[35] , \R_DATA_TEMPR13[34] }), 
        .B_DOUT({nc7352, nc7353, nc7354, nc7355, nc7356, nc7357, 
        nc7358, nc7359, nc7360, nc7361, nc7362, nc7363, nc7364, nc7365, 
        nc7366, nc7367, nc7368, nc7369, nc7370, nc7371}), .DB_DETECT(
        \DB_DETECT[13][17] ), .SB_CORRECT(\SB_CORRECT[13][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_30 (.A(\R_DATA_TEMPR8[14] ), .B(\R_DATA_TEMPR9[14] ), .C(
        \R_DATA_TEMPR10[14] ), .D(\R_DATA_TEMPR11[14] ), .Y(OR4_30_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C7 (.A_DOUT({nc7372, 
        nc7373, nc7374, nc7375, nc7376, nc7377, nc7378, nc7379, nc7380, 
        nc7381, nc7382, nc7383, nc7384, nc7385, nc7386, nc7387, nc7388, 
        nc7389, \R_DATA_TEMPR2[15] , \R_DATA_TEMPR2[14] }), .B_DOUT({
        nc7390, nc7391, nc7392, nc7393, nc7394, nc7395, nc7396, nc7397, 
        nc7398, nc7399, nc7400, nc7401, nc7402, nc7403, nc7404, nc7405, 
        nc7406, nc7407, nc7408, nc7409}), .DB_DETECT(\DB_DETECT[2][7] )
        , .SB_CORRECT(\SB_CORRECT[2][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_297 (.A(OR4_287_Y), .B(OR4_283_Y), .C(OR4_255_Y), .D(
        OR4_353_Y), .Y(OR4_297_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C19 (.A_DOUT({nc7410, 
        nc7411, nc7412, nc7413, nc7414, nc7415, nc7416, nc7417, nc7418, 
        nc7419, nc7420, nc7421, nc7422, nc7423, nc7424, nc7425, nc7426, 
        nc7427, \R_DATA_TEMPR3[39] , \R_DATA_TEMPR3[38] }), .B_DOUT({
        nc7428, nc7429, nc7430, nc7431, nc7432, nc7433, nc7434, nc7435, 
        nc7436, nc7437, nc7438, nc7439, nc7440, nc7441, nc7442, nc7443, 
        nc7444, nc7445, nc7446, nc7447}), .DB_DETECT(
        \DB_DETECT[3][19] ), .SB_CORRECT(\SB_CORRECT[3][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_37 (.A(\R_DATA_TEMPR12[20] ), .B(\R_DATA_TEMPR13[20] ), .C(
        \R_DATA_TEMPR14[20] ), .D(\R_DATA_TEMPR15[20] ), .Y(OR4_37_Y));
    OR4 OR4_197 (.A(\R_DATA_TEMPR8[9] ), .B(\R_DATA_TEMPR9[9] ), .C(
        \R_DATA_TEMPR10[9] ), .D(\R_DATA_TEMPR11[9] ), .Y(OR4_197_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C9 (.A_DOUT({nc7448, 
        nc7449, nc7450, nc7451, nc7452, nc7453, nc7454, nc7455, nc7456, 
        nc7457, nc7458, nc7459, nc7460, nc7461, nc7462, nc7463, nc7464, 
        nc7465, \R_DATA_TEMPR13[19] , \R_DATA_TEMPR13[18] }), .B_DOUT({
        nc7466, nc7467, nc7468, nc7469, nc7470, nc7471, nc7472, nc7473, 
        nc7474, nc7475, nc7476, nc7477, nc7478, nc7479, nc7480, nc7481, 
        nc7482, nc7483, nc7484, nc7485}), .DB_DETECT(
        \DB_DETECT[13][9] ), .SB_CORRECT(\SB_CORRECT[13][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_357 (.A(\R_DATA_TEMPR4[33] ), .B(\R_DATA_TEMPR5[33] ), .C(
        \R_DATA_TEMPR6[33] ), .D(\R_DATA_TEMPR7[33] ), .Y(OR4_357_Y));
    OR4 OR4_150 (.A(\R_DATA_TEMPR4[18] ), .B(\R_DATA_TEMPR5[18] ), .C(
        \R_DATA_TEMPR6[18] ), .D(\R_DATA_TEMPR7[18] ), .Y(OR4_150_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[5]  (.A(CFG2_6_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[5] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C12 (.A_DOUT({nc7486, 
        nc7487, nc7488, nc7489, nc7490, nc7491, nc7492, nc7493, nc7494, 
        nc7495, nc7496, nc7497, nc7498, nc7499, nc7500, nc7501, nc7502, 
        nc7503, \R_DATA_TEMPR0[25] , \R_DATA_TEMPR0[24] }), .B_DOUT({
        nc7504, nc7505, nc7506, nc7507, nc7508, nc7509, nc7510, nc7511, 
        nc7512, nc7513, nc7514, nc7515, nc7516, nc7517, nc7518, nc7519, 
        nc7520, nc7521, nc7522, nc7523}), .DB_DETECT(
        \DB_DETECT[0][12] ), .SB_CORRECT(\SB_CORRECT[0][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h2) )  CFG2_7 (.A(W_ADDR[16]), .B(W_ADDR[15]), .Y(
        CFG2_7_Y));
    OR4 OR4_163 (.A(\R_DATA_TEMPR24[22] ), .B(\R_DATA_TEMPR25[22] ), 
        .C(\R_DATA_TEMPR26[22] ), .D(\R_DATA_TEMPR27[22] ), .Y(
        OR4_163_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C4 (.A_DOUT({nc7524, 
        nc7525, nc7526, nc7527, nc7528, nc7529, nc7530, nc7531, nc7532, 
        nc7533, nc7534, nc7535, nc7536, nc7537, nc7538, nc7539, nc7540, 
        nc7541, \R_DATA_TEMPR2[9] , \R_DATA_TEMPR2[8] }), .B_DOUT({
        nc7542, nc7543, nc7544, nc7545, nc7546, nc7547, nc7548, nc7549, 
        nc7550, nc7551, nc7552, nc7553, nc7554, nc7555, nc7556, nc7557, 
        nc7558, nc7559, nc7560, nc7561}), .DB_DETECT(\DB_DETECT[2][4] )
        , .SB_CORRECT(\SB_CORRECT[2][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_343 (.A(OR4_50_Y), .B(OR2_5_Y), .C(\R_DATA_TEMPR22[5] ), 
        .D(\R_DATA_TEMPR23[5] ), .Y(OR4_343_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[7]  (.A(CFG2_5_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[7] ));
    OR4 OR4_336 (.A(\R_DATA_TEMPR0[13] ), .B(\R_DATA_TEMPR1[13] ), .C(
        \R_DATA_TEMPR2[13] ), .D(\R_DATA_TEMPR3[13] ), .Y(OR4_336_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C3 (.A_DOUT({nc7562, 
        nc7563, nc7564, nc7565, nc7566, nc7567, nc7568, nc7569, nc7570, 
        nc7571, nc7572, nc7573, nc7574, nc7575, nc7576, nc7577, nc7578, 
        nc7579, \R_DATA_TEMPR6[7] , \R_DATA_TEMPR6[6] }), .B_DOUT({
        nc7580, nc7581, nc7582, nc7583, nc7584, nc7585, nc7586, nc7587, 
        nc7588, nc7589, nc7590, nc7591, nc7592, nc7593, nc7594, nc7595, 
        nc7596, nc7597, nc7598, nc7599}), .DB_DETECT(\DB_DETECT[6][3] )
        , .SB_CORRECT(\SB_CORRECT[6][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_294 (.A(OR4_266_Y), .B(OR4_186_Y), .C(OR4_270_Y), .D(
        OR4_73_Y), .Y(OR4_294_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C2 (.A_DOUT({nc7600, 
        nc7601, nc7602, nc7603, nc7604, nc7605, nc7606, nc7607, nc7608, 
        nc7609, nc7610, nc7611, nc7612, nc7613, nc7614, nc7615, nc7616, 
        nc7617, \R_DATA_TEMPR14[5] , \R_DATA_TEMPR14[4] }), .B_DOUT({
        nc7618, nc7619, nc7620, nc7621, nc7622, nc7623, nc7624, nc7625, 
        nc7626, nc7627, nc7628, nc7629, nc7630, nc7631, nc7632, nc7633, 
        nc7634, nc7635, nc7636, nc7637}), .DB_DETECT(
        \DB_DETECT[14][2] ), .SB_CORRECT(\SB_CORRECT[14][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[24]  (.A(OR4_308_Y), .B(OR4_181_Y), .C(OR4_1_Y), 
        .D(OR4_152_Y), .Y(R_DATA[24]));
    OR4 OR4_85 (.A(\R_DATA_TEMPR12[28] ), .B(\R_DATA_TEMPR13[28] ), .C(
        \R_DATA_TEMPR14[28] ), .D(\R_DATA_TEMPR15[28] ), .Y(OR4_85_Y));
    OR4 OR4_146 (.A(\R_DATA_TEMPR4[21] ), .B(\R_DATA_TEMPR5[21] ), .C(
        \R_DATA_TEMPR6[21] ), .D(\R_DATA_TEMPR7[21] ), .Y(OR4_146_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C4 (.A_DOUT({nc7638, 
        nc7639, nc7640, nc7641, nc7642, nc7643, nc7644, nc7645, nc7646, 
        nc7647, nc7648, nc7649, nc7650, nc7651, nc7652, nc7653, nc7654, 
        nc7655, \R_DATA_TEMPR19[9] , \R_DATA_TEMPR19[8] }), .B_DOUT({
        nc7656, nc7657, nc7658, nc7659, nc7660, nc7661, nc7662, nc7663, 
        nc7664, nc7665, nc7666, nc7667, nc7668, nc7669, nc7670, nc7671, 
        nc7672, nc7673, nc7674, nc7675}), .DB_DETECT(
        \DB_DETECT[19][4] ), .SB_CORRECT(\SB_CORRECT[19][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_158 (.A(\R_DATA_TEMPR4[6] ), .B(\R_DATA_TEMPR5[6] ), .C(
        \R_DATA_TEMPR6[6] ), .D(\R_DATA_TEMPR7[6] ), .Y(OR4_158_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_256_Y), .B(OR4_245_Y), .C(OR4_196_Y), 
        .D(OR4_29_Y), .Y(R_DATA[12]));
    OR4 OR4_69 (.A(\R_DATA_TEMPR16[6] ), .B(\R_DATA_TEMPR17[6] ), .C(
        \R_DATA_TEMPR18[6] ), .D(\R_DATA_TEMPR19[6] ), .Y(OR4_69_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C2 (.A_DOUT({nc7676, 
        nc7677, nc7678, nc7679, nc7680, nc7681, nc7682, nc7683, nc7684, 
        nc7685, nc7686, nc7687, nc7688, nc7689, nc7690, nc7691, nc7692, 
        nc7693, \R_DATA_TEMPR23[5] , \R_DATA_TEMPR23[4] }), .B_DOUT({
        nc7694, nc7695, nc7696, nc7697, nc7698, nc7699, nc7700, nc7701, 
        nc7702, nc7703, nc7704, nc7705, nc7706, nc7707, nc7708, nc7709, 
        nc7710, nc7711, nc7712, nc7713}), .DB_DETECT(
        \DB_DETECT[23][2] ), .SB_CORRECT(\SB_CORRECT[23][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_227 (.A(\R_DATA_TEMPR8[23] ), .B(\R_DATA_TEMPR9[23] ), .C(
        \R_DATA_TEMPR10[23] ), .D(\R_DATA_TEMPR11[23] ), .Y(OR4_227_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C9 (.A_DOUT({nc7714, 
        nc7715, nc7716, nc7717, nc7718, nc7719, nc7720, nc7721, nc7722, 
        nc7723, nc7724, nc7725, nc7726, nc7727, nc7728, nc7729, nc7730, 
        nc7731, \R_DATA_TEMPR30[19] , \R_DATA_TEMPR30[18] }), .B_DOUT({
        nc7732, nc7733, nc7734, nc7735, nc7736, nc7737, nc7738, nc7739, 
        nc7740, nc7741, nc7742, nc7743, nc7744, nc7745, nc7746, nc7747, 
        nc7748, nc7749, nc7750, nc7751}), .DB_DETECT(
        \DB_DETECT[30][9] ), .SB_CORRECT(\SB_CORRECT[30][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][9] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_127 (.A(\R_DATA_TEMPR0[11] ), .B(\R_DATA_TEMPR1[11] ), .C(
        \R_DATA_TEMPR2[11] ), .D(\R_DATA_TEMPR3[11] ), .Y(OR4_127_Y));
    OR4 OR4_348 (.A(\R_DATA_TEMPR8[33] ), .B(\R_DATA_TEMPR9[33] ), .C(
        \R_DATA_TEMPR10[33] ), .D(\R_DATA_TEMPR11[33] ), .Y(OR4_348_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C6 (.A_DOUT({nc7752, 
        nc7753, nc7754, nc7755, nc7756, nc7757, nc7758, nc7759, nc7760, 
        nc7761, nc7762, nc7763, nc7764, nc7765, nc7766, nc7767, nc7768, 
        nc7769, \R_DATA_TEMPR11[13] , \R_DATA_TEMPR11[12] }), .B_DOUT({
        nc7770, nc7771, nc7772, nc7773, nc7774, nc7775, nc7776, nc7777, 
        nc7778, nc7779, nc7780, nc7781, nc7782, nc7783, nc7784, nc7785, 
        nc7786, nc7787, nc7788, nc7789}), .DB_DETECT(
        \DB_DETECT[11][6] ), .SB_CORRECT(\SB_CORRECT[11][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C4 (.A_DOUT({nc7790, 
        nc7791, nc7792, nc7793, nc7794, nc7795, nc7796, nc7797, nc7798, 
        nc7799, nc7800, nc7801, nc7802, nc7803, nc7804, nc7805, nc7806, 
        nc7807, \R_DATA_TEMPR25[9] , \R_DATA_TEMPR25[8] }), .B_DOUT({
        nc7808, nc7809, nc7810, nc7811, nc7812, nc7813, nc7814, nc7815, 
        nc7816, nc7817, nc7818, nc7819, nc7820, nc7821, nc7822, nc7823, 
        nc7824, nc7825, nc7826, nc7827}), .DB_DETECT(
        \DB_DETECT[25][4] ), .SB_CORRECT(\SB_CORRECT[25][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_162 (.A(\R_DATA_TEMPR28[36] ), .B(\R_DATA_TEMPR29[36] ), 
        .C(\R_DATA_TEMPR30[36] ), .D(\R_DATA_TEMPR31[36] ), .Y(
        OR4_162_Y));
    OR4 OR4_282 (.A(\R_DATA_TEMPR24[32] ), .B(\R_DATA_TEMPR25[32] ), 
        .C(\R_DATA_TEMPR26[32] ), .D(\R_DATA_TEMPR27[32] ), .Y(
        OR4_282_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C19 (.A_DOUT({
        nc7828, nc7829, nc7830, nc7831, nc7832, nc7833, nc7834, nc7835, 
        nc7836, nc7837, nc7838, nc7839, nc7840, nc7841, nc7842, nc7843, 
        nc7844, nc7845, \R_DATA_TEMPR26[39] , \R_DATA_TEMPR26[38] }), 
        .B_DOUT({nc7846, nc7847, nc7848, nc7849, nc7850, nc7851, 
        nc7852, nc7853, nc7854, nc7855, nc7856, nc7857, nc7858, nc7859, 
        nc7860, nc7861, nc7862, nc7863, nc7864, nc7865}), .DB_DETECT(
        \DB_DETECT[26][19] ), .SB_CORRECT(\SB_CORRECT[26][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_316 (.A(\R_DATA_TEMPR8[3] ), .B(\R_DATA_TEMPR9[3] ), .C(
        \R_DATA_TEMPR10[3] ), .D(\R_DATA_TEMPR11[3] ), .Y(OR4_316_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C6 (.A_DOUT({nc7866, 
        nc7867, nc7868, nc7869, nc7870, nc7871, nc7872, nc7873, nc7874, 
        nc7875, nc7876, nc7877, nc7878, nc7879, nc7880, nc7881, nc7882, 
        nc7883, \R_DATA_TEMPR17[13] , \R_DATA_TEMPR17[12] }), .B_DOUT({
        nc7884, nc7885, nc7886, nc7887, nc7888, nc7889, nc7890, nc7891, 
        nc7892, nc7893, nc7894, nc7895, nc7896, nc7897, nc7898, nc7899, 
        nc7900, nc7901, nc7902, nc7903}), .DB_DETECT(
        \DB_DETECT[17][6] ), .SB_CORRECT(\SB_CORRECT[17][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C18 (.A_DOUT({
        nc7904, nc7905, nc7906, nc7907, nc7908, nc7909, nc7910, nc7911, 
        nc7912, nc7913, nc7914, nc7915, nc7916, nc7917, nc7918, nc7919, 
        nc7920, nc7921, \R_DATA_TEMPR11[37] , \R_DATA_TEMPR11[36] }), 
        .B_DOUT({nc7922, nc7923, nc7924, nc7925, nc7926, nc7927, 
        nc7928, nc7929, nc7930, nc7931, nc7932, nc7933, nc7934, nc7935, 
        nc7936, nc7937, nc7938, nc7939, nc7940, nc7941}), .DB_DETECT(
        \DB_DETECT[11][18] ), .SB_CORRECT(\SB_CORRECT[11][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_134 (.A(\R_DATA_TEMPR24[8] ), .B(\R_DATA_TEMPR25[8] ), .C(
        \R_DATA_TEMPR26[8] ), .D(\R_DATA_TEMPR27[8] ), .Y(OR4_134_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C6 (.A_DOUT({nc7942, 
        nc7943, nc7944, nc7945, nc7946, nc7947, nc7948, nc7949, nc7950, 
        nc7951, nc7952, nc7953, nc7954, nc7955, nc7956, nc7957, nc7958, 
        nc7959, \R_DATA_TEMPR30[13] , \R_DATA_TEMPR30[12] }), .B_DOUT({
        nc7960, nc7961, nc7962, nc7963, nc7964, nc7965, nc7966, nc7967, 
        nc7968, nc7969, nc7970, nc7971, nc7972, nc7973, nc7974, nc7975, 
        nc7976, nc7977, nc7978, nc7979}), .DB_DETECT(
        \DB_DETECT[30][6] ), .SB_CORRECT(\SB_CORRECT[30][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_35 (.A(\R_DATA_TEMPR20[0] ), .B(\R_DATA_TEMPR21[0] ), .Y(
        OR2_35_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C17 (.A_DOUT({
        nc7980, nc7981, nc7982, nc7983, nc7984, nc7985, nc7986, nc7987, 
        nc7988, nc7989, nc7990, nc7991, nc7992, nc7993, nc7994, nc7995, 
        nc7996, nc7997, \R_DATA_TEMPR10[35] , \R_DATA_TEMPR10[34] }), 
        .B_DOUT({nc7998, nc7999, nc8000, nc8001, nc8002, nc8003, 
        nc8004, nc8005, nc8006, nc8007, nc8008, nc8009, nc8010, nc8011, 
        nc8012, nc8013, nc8014, nc8015, nc8016, nc8017}), .DB_DETECT(
        \DB_DETECT[10][17] ), .SB_CORRECT(\SB_CORRECT[10][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C14 (.A_DOUT({nc8018, 
        nc8019, nc8020, nc8021, nc8022, nc8023, nc8024, nc8025, nc8026, 
        nc8027, nc8028, nc8029, nc8030, nc8031, nc8032, nc8033, nc8034, 
        nc8035, \R_DATA_TEMPR2[29] , \R_DATA_TEMPR2[28] }), .B_DOUT({
        nc8036, nc8037, nc8038, nc8039, nc8040, nc8041, nc8042, nc8043, 
        nc8044, nc8045, nc8046, nc8047, nc8048, nc8049, nc8050, nc8051, 
        nc8052, nc8053, nc8054, nc8055}), .DB_DETECT(
        \DB_DETECT[2][14] ), .SB_CORRECT(\SB_CORRECT[2][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_103 (.A(OR4_144_Y), .B(OR2_11_Y), .C(\R_DATA_TEMPR22[30] ), 
        .D(\R_DATA_TEMPR23[30] ), .Y(OR4_103_Y));
    OR4 OR4_224 (.A(\R_DATA_TEMPR24[7] ), .B(\R_DATA_TEMPR25[7] ), .C(
        \R_DATA_TEMPR26[7] ), .D(\R_DATA_TEMPR27[7] ), .Y(OR4_224_Y));
    OR4 OR4_149 (.A(\R_DATA_TEMPR28[4] ), .B(\R_DATA_TEMPR29[4] ), .C(
        \R_DATA_TEMPR30[4] ), .D(\R_DATA_TEMPR31[4] ), .Y(OR4_149_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C14 (.A_DOUT({
        nc8056, nc8057, nc8058, nc8059, nc8060, nc8061, nc8062, nc8063, 
        nc8064, nc8065, nc8066, nc8067, nc8068, nc8069, nc8070, nc8071, 
        nc8072, nc8073, \R_DATA_TEMPR17[29] , \R_DATA_TEMPR17[28] }), 
        .B_DOUT({nc8074, nc8075, nc8076, nc8077, nc8078, nc8079, 
        nc8080, nc8081, nc8082, nc8083, nc8084, nc8085, nc8086, nc8087, 
        nc8088, nc8089, nc8090, nc8091, nc8092, nc8093}), .DB_DETECT(
        \DB_DETECT[17][14] ), .SB_CORRECT(\SB_CORRECT[17][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[13]  (.A(OR4_212_Y), .B(OR4_130_Y), .C(OR4_114_Y), 
        .D(OR4_106_Y), .Y(R_DATA[13]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0 (.A_DOUT({nc8094, 
        nc8095, nc8096, nc8097, nc8098, nc8099, nc8100, nc8101, nc8102, 
        nc8103, nc8104, nc8105, nc8106, nc8107, nc8108, nc8109, nc8110, 
        nc8111, \R_DATA_TEMPR25[1] , \R_DATA_TEMPR25[0] }), .B_DOUT({
        nc8112, nc8113, nc8114, nc8115, nc8116, nc8117, nc8118, nc8119, 
        nc8120, nc8121, nc8122, nc8123, nc8124, nc8125, nc8126, nc8127, 
        nc8128, nc8129, nc8130, nc8131}), .DB_DETECT(
        \DB_DETECT[25][0] ), .SB_CORRECT(\SB_CORRECT[25][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][0] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_173 (.A(\R_DATA_TEMPR28[18] ), .B(\R_DATA_TEMPR29[18] ), 
        .C(\R_DATA_TEMPR30[18] ), .D(\R_DATA_TEMPR31[18] ), .Y(
        OR4_173_Y));
    OR4 OR4_269 (.A(\R_DATA_TEMPR28[8] ), .B(\R_DATA_TEMPR29[8] ), .C(
        \R_DATA_TEMPR30[8] ), .D(\R_DATA_TEMPR31[8] ), .Y(OR4_269_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C2 (.A_DOUT({nc8132, 
        nc8133, nc8134, nc8135, nc8136, nc8137, nc8138, nc8139, nc8140, 
        nc8141, nc8142, nc8143, nc8144, nc8145, nc8146, nc8147, nc8148, 
        nc8149, \R_DATA_TEMPR3[5] , \R_DATA_TEMPR3[4] }), .B_DOUT({
        nc8150, nc8151, nc8152, nc8153, nc8154, nc8155, nc8156, nc8157, 
        nc8158, nc8159, nc8160, nc8161, nc8162, nc8163, nc8164, nc8165, 
        nc8166, nc8167, nc8168, nc8169}), .DB_DETECT(\DB_DETECT[3][2] )
        , .SB_CORRECT(\SB_CORRECT[3][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1 (.A_DOUT({nc8170, 
        nc8171, nc8172, nc8173, nc8174, nc8175, nc8176, nc8177, nc8178, 
        nc8179, nc8180, nc8181, nc8182, nc8183, nc8184, nc8185, nc8186, 
        nc8187, \R_DATA_TEMPR4[3] , \R_DATA_TEMPR4[2] }), .B_DOUT({
        nc8188, nc8189, nc8190, nc8191, nc8192, nc8193, nc8194, nc8195, 
        nc8196, nc8197, nc8198, nc8199, nc8200, nc8201, nc8202, nc8203, 
        nc8204, nc8205, nc8206, nc8207}), .DB_DETECT(\DB_DETECT[4][1] )
        , .SB_CORRECT(\SB_CORRECT[4][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_62 (.A(\R_DATA_TEMPR16[22] ), .B(\R_DATA_TEMPR17[22] ), .C(
        \R_DATA_TEMPR18[22] ), .D(\R_DATA_TEMPR19[22] ), .Y(OR4_62_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C10 (.A_DOUT({
        nc8208, nc8209, nc8210, nc8211, nc8212, nc8213, nc8214, nc8215, 
        nc8216, nc8217, nc8218, nc8219, nc8220, nc8221, nc8222, nc8223, 
        nc8224, nc8225, \R_DATA_TEMPR18[21] , \R_DATA_TEMPR18[20] }), 
        .B_DOUT({nc8226, nc8227, nc8228, nc8229, nc8230, nc8231, 
        nc8232, nc8233, nc8234, nc8235, nc8236, nc8237, nc8238, nc8239, 
        nc8240, nc8241, nc8242, nc8243, nc8244, nc8245}), .DB_DETECT(
        \DB_DETECT[18][10] ), .SB_CORRECT(\SB_CORRECT[18][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C8 (.A_DOUT({nc8246, 
        nc8247, nc8248, nc8249, nc8250, nc8251, nc8252, nc8253, nc8254, 
        nc8255, nc8256, nc8257, nc8258, nc8259, nc8260, nc8261, nc8262, 
        nc8263, \R_DATA_TEMPR29[17] , \R_DATA_TEMPR29[16] }), .B_DOUT({
        nc8264, nc8265, nc8266, nc8267, nc8268, nc8269, nc8270, nc8271, 
        nc8272, nc8273, nc8274, nc8275, nc8276, nc8277, nc8278, nc8279, 
        nc8280, nc8281, nc8282, nc8283}), .DB_DETECT(
        \DB_DETECT[29][8] ), .SB_CORRECT(\SB_CORRECT[29][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_38 (.A(\R_DATA_TEMPR12[39] ), .B(\R_DATA_TEMPR13[39] ), .C(
        \R_DATA_TEMPR14[39] ), .D(\R_DATA_TEMPR15[39] ), .Y(OR4_38_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C3 (.A_DOUT({nc8284, 
        nc8285, nc8286, nc8287, nc8288, nc8289, nc8290, nc8291, nc8292, 
        nc8293, nc8294, nc8295, nc8296, nc8297, nc8298, nc8299, nc8300, 
        nc8301, \R_DATA_TEMPR18[7] , \R_DATA_TEMPR18[6] }), .B_DOUT({
        nc8302, nc8303, nc8304, nc8305, nc8306, nc8307, nc8308, nc8309, 
        nc8310, nc8311, nc8312, nc8313, nc8314, nc8315, nc8316, nc8317, 
        nc8318, nc8319, nc8320, nc8321}), .DB_DETECT(
        \DB_DETECT[18][3] ), .SB_CORRECT(\SB_CORRECT[18][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C15 (.A_DOUT({
        nc8322, nc8323, nc8324, nc8325, nc8326, nc8327, nc8328, nc8329, 
        nc8330, nc8331, nc8332, nc8333, nc8334, nc8335, nc8336, nc8337, 
        nc8338, nc8339, \R_DATA_TEMPR18[31] , \R_DATA_TEMPR18[30] }), 
        .B_DOUT({nc8340, nc8341, nc8342, nc8343, nc8344, nc8345, 
        nc8346, nc8347, nc8348, nc8349, nc8350, nc8351, nc8352, nc8353, 
        nc8354, nc8355, nc8356, nc8357, nc8358, nc8359}), .DB_DETECT(
        \DB_DETECT[18][15] ), .SB_CORRECT(\SB_CORRECT[18][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][15] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_325 (.A(OR4_101_Y), .B(OR2_25_Y), .C(\R_DATA_TEMPR22[7] ), 
        .D(\R_DATA_TEMPR23[7] ), .Y(OR4_325_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C11 (.A_DOUT({
        nc8360, nc8361, nc8362, nc8363, nc8364, nc8365, nc8366, nc8367, 
        nc8368, nc8369, nc8370, nc8371, nc8372, nc8373, nc8374, nc8375, 
        nc8376, nc8377, \R_DATA_TEMPR19[23] , \R_DATA_TEMPR19[22] }), 
        .B_DOUT({nc8378, nc8379, nc8380, nc8381, nc8382, nc8383, 
        nc8384, nc8385, nc8386, nc8387, nc8388, nc8389, nc8390, nc8391, 
        nc8392, nc8393, nc8394, nc8395, nc8396, nc8397}), .DB_DETECT(
        \DB_DETECT[19][11] ), .SB_CORRECT(\SB_CORRECT[19][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C14 (.A_DOUT({nc8398, 
        nc8399, nc8400, nc8401, nc8402, nc8403, nc8404, nc8405, nc8406, 
        nc8407, nc8408, nc8409, nc8410, nc8411, nc8412, nc8413, nc8414, 
        nc8415, \R_DATA_TEMPR7[29] , \R_DATA_TEMPR7[28] }), .B_DOUT({
        nc8416, nc8417, nc8418, nc8419, nc8420, nc8421, nc8422, nc8423, 
        nc8424, nc8425, nc8426, nc8427, nc8428, nc8429, nc8430, nc8431, 
        nc8432, nc8433, nc8434, nc8435}), .DB_DETECT(
        \DB_DETECT[7][14] ), .SB_CORRECT(\SB_CORRECT[7][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C18 (.A_DOUT({
        nc8436, nc8437, nc8438, nc8439, nc8440, nc8441, nc8442, nc8443, 
        nc8444, nc8445, nc8446, nc8447, nc8448, nc8449, nc8450, nc8451, 
        nc8452, nc8453, \R_DATA_TEMPR26[37] , \R_DATA_TEMPR26[36] }), 
        .B_DOUT({nc8454, nc8455, nc8456, nc8457, nc8458, nc8459, 
        nc8460, nc8461, nc8462, nc8463, nc8464, nc8465, nc8466, nc8467, 
        nc8468, nc8469, nc8470, nc8471, nc8472, nc8473}), .DB_DETECT(
        \DB_DETECT[26][18] ), .SB_CORRECT(\SB_CORRECT[26][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C12 (.A_DOUT({
        nc8474, nc8475, nc8476, nc8477, nc8478, nc8479, nc8480, nc8481, 
        nc8482, nc8483, nc8484, nc8485, nc8486, nc8487, nc8488, nc8489, 
        nc8490, nc8491, \R_DATA_TEMPR13[25] , \R_DATA_TEMPR13[24] }), 
        .B_DOUT({nc8492, nc8493, nc8494, nc8495, nc8496, nc8497, 
        nc8498, nc8499, nc8500, nc8501, nc8502, nc8503, nc8504, nc8505, 
        nc8506, nc8507, nc8508, nc8509, nc8510, nc8511}), .DB_DETECT(
        \DB_DETECT[13][12] ), .SB_CORRECT(\SB_CORRECT[13][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1 (.A_DOUT({nc8512, 
        nc8513, nc8514, nc8515, nc8516, nc8517, nc8518, nc8519, nc8520, 
        nc8521, nc8522, nc8523, nc8524, nc8525, nc8526, nc8527, nc8528, 
        nc8529, \R_DATA_TEMPR11[3] , \R_DATA_TEMPR11[2] }), .B_DOUT({
        nc8530, nc8531, nc8532, nc8533, nc8534, nc8535, nc8536, nc8537, 
        nc8538, nc8539, nc8540, nc8541, nc8542, nc8543, nc8544, nc8545, 
        nc8546, nc8547, nc8548, nc8549}), .DB_DETECT(
        \DB_DETECT[11][1] ), .SB_CORRECT(\SB_CORRECT[11][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][1] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C11 (.A_DOUT({
        nc8550, nc8551, nc8552, nc8553, nc8554, nc8555, nc8556, nc8557, 
        nc8558, nc8559, nc8560, nc8561, nc8562, nc8563, nc8564, nc8565, 
        nc8566, nc8567, \R_DATA_TEMPR23[23] , \R_DATA_TEMPR23[22] }), 
        .B_DOUT({nc8568, nc8569, nc8570, nc8571, nc8572, nc8573, 
        nc8574, nc8575, nc8576, nc8577, nc8578, nc8579, nc8580, nc8581, 
        nc8582, nc8583, nc8584, nc8585, nc8586, nc8587}), .DB_DETECT(
        \DB_DETECT[23][11] ), .SB_CORRECT(\SB_CORRECT[23][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C3 (.A_DOUT({nc8588, 
        nc8589, nc8590, nc8591, nc8592, nc8593, nc8594, nc8595, nc8596, 
        nc8597, nc8598, nc8599, nc8600, nc8601, nc8602, nc8603, nc8604, 
        nc8605, \R_DATA_TEMPR31[7] , \R_DATA_TEMPR31[6] }), .B_DOUT({
        nc8606, nc8607, nc8608, nc8609, nc8610, nc8611, nc8612, nc8613, 
        nc8614, nc8615, nc8616, nc8617, nc8618, nc8619, nc8620, nc8621, 
        nc8622, nc8623, nc8624, nc8625}), .DB_DETECT(
        \DB_DETECT[31][3] ), .SB_CORRECT(\SB_CORRECT[31][3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][3] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_114 (.A(\R_DATA_TEMPR24[13] ), .B(\R_DATA_TEMPR25[13] ), 
        .C(\R_DATA_TEMPR26[13] ), .D(\R_DATA_TEMPR27[13] ), .Y(
        OR4_114_Y));
    OR4 OR4_155 (.A(\R_DATA_TEMPR16[29] ), .B(\R_DATA_TEMPR17[29] ), 
        .C(\R_DATA_TEMPR18[29] ), .D(\R_DATA_TEMPR19[29] ), .Y(
        OR4_155_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C8 (.A_DOUT({nc8626, 
        nc8627, nc8628, nc8629, nc8630, nc8631, nc8632, nc8633, nc8634, 
        nc8635, nc8636, nc8637, nc8638, nc8639, nc8640, nc8641, nc8642, 
        nc8643, \R_DATA_TEMPR10[17] , \R_DATA_TEMPR10[16] }), .B_DOUT({
        nc8644, nc8645, nc8646, nc8647, nc8648, nc8649, nc8650, nc8651, 
        nc8652, nc8653, nc8654, nc8655, nc8656, nc8657, nc8658, nc8659, 
        nc8660, nc8661, nc8662, nc8663}), .DB_DETECT(
        \DB_DETECT[10][8] ), .SB_CORRECT(\SB_CORRECT[10][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C17 (.A_DOUT({nc8664, 
        nc8665, nc8666, nc8667, nc8668, nc8669, nc8670, nc8671, nc8672, 
        nc8673, nc8674, nc8675, nc8676, nc8677, nc8678, nc8679, nc8680, 
        nc8681, \R_DATA_TEMPR4[35] , \R_DATA_TEMPR4[34] }), .B_DOUT({
        nc8682, nc8683, nc8684, nc8685, nc8686, nc8687, nc8688, nc8689, 
        nc8690, nc8691, nc8692, nc8693, nc8694, nc8695, nc8696, nc8697, 
        nc8698, nc8699, nc8700, nc8701}), .DB_DETECT(
        \DB_DETECT[4][17] ), .SB_CORRECT(\SB_CORRECT[4][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C4 (.A_DOUT({nc8702, 
        nc8703, nc8704, nc8705, nc8706, nc8707, nc8708, nc8709, nc8710, 
        nc8711, nc8712, nc8713, nc8714, nc8715, nc8716, nc8717, nc8718, 
        nc8719, \R_DATA_TEMPR22[9] , \R_DATA_TEMPR22[8] }), .B_DOUT({
        nc8720, nc8721, nc8722, nc8723, nc8724, nc8725, nc8726, nc8727, 
        nc8728, nc8729, nc8730, nc8731, nc8732, nc8733, nc8734, nc8735, 
        nc8736, nc8737, nc8738, nc8739}), .DB_DETECT(
        \DB_DETECT[22][4] ), .SB_CORRECT(\SB_CORRECT[22][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C11 (.A_DOUT({nc8740, 
        nc8741, nc8742, nc8743, nc8744, nc8745, nc8746, nc8747, nc8748, 
        nc8749, nc8750, nc8751, nc8752, nc8753, nc8754, nc8755, nc8756, 
        nc8757, \R_DATA_TEMPR9[23] , \R_DATA_TEMPR9[22] }), .B_DOUT({
        nc8758, nc8759, nc8760, nc8761, nc8762, nc8763, nc8764, nc8765, 
        nc8766, nc8767, nc8768, nc8769, nc8770, nc8771, nc8772, nc8773, 
        nc8774, nc8775, nc8776, nc8777}), .DB_DETECT(
        \DB_DETECT[9][11] ), .SB_CORRECT(\SB_CORRECT[9][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C2 (.A_DOUT({nc8778, 
        nc8779, nc8780, nc8781, nc8782, nc8783, nc8784, nc8785, nc8786, 
        nc8787, nc8788, nc8789, nc8790, nc8791, nc8792, nc8793, nc8794, 
        nc8795, \R_DATA_TEMPR22[5] , \R_DATA_TEMPR22[4] }), .B_DOUT({
        nc8796, nc8797, nc8798, nc8799, nc8800, nc8801, nc8802, nc8803, 
        nc8804, nc8805, nc8806, nc8807, nc8808, nc8809, nc8810, nc8811, 
        nc8812, nc8813, nc8814, nc8815}), .DB_DETECT(
        \DB_DETECT[22][2] ), .SB_CORRECT(\SB_CORRECT[22][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C16 (.A_DOUT({nc8816, 
        nc8817, nc8818, nc8819, nc8820, nc8821, nc8822, nc8823, nc8824, 
        nc8825, nc8826, nc8827, nc8828, nc8829, nc8830, nc8831, nc8832, 
        nc8833, \R_DATA_TEMPR1[33] , \R_DATA_TEMPR1[32] }), .B_DOUT({
        nc8834, nc8835, nc8836, nc8837, nc8838, nc8839, nc8840, nc8841, 
        nc8842, nc8843, nc8844, nc8845, nc8846, nc8847, nc8848, nc8849, 
        nc8850, nc8851, nc8852, nc8853}), .DB_DETECT(
        \DB_DETECT[1][16] ), .SB_CORRECT(\SB_CORRECT[1][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_102 (.A(\R_DATA_TEMPR8[18] ), .B(\R_DATA_TEMPR9[18] ), .C(
        \R_DATA_TEMPR10[18] ), .D(\R_DATA_TEMPR11[18] ), .Y(OR4_102_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C19 (.A_DOUT({nc8854, 
        nc8855, nc8856, nc8857, nc8858, nc8859, nc8860, nc8861, nc8862, 
        nc8863, nc8864, nc8865, nc8866, nc8867, nc8868, nc8869, nc8870, 
        nc8871, \R_DATA_TEMPR0[39] , \R_DATA_TEMPR0[38] }), .B_DOUT({
        nc8872, nc8873, nc8874, nc8875, nc8876, nc8877, nc8878, nc8879, 
        nc8880, nc8881, nc8882, nc8883, nc8884, nc8885, nc8886, nc8887, 
        nc8888, nc8889, nc8890, nc8891}), .DB_DETECT(
        \DB_DETECT[0][19] ), .SB_CORRECT(\SB_CORRECT[0][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    INV \INVBLKY0[0]  (.A(R_ADDR[13]), .Y(\BLKY0[0] ));
    OR4 OR4_172 (.A(\R_DATA_TEMPR16[32] ), .B(\R_DATA_TEMPR17[32] ), 
        .C(\R_DATA_TEMPR18[32] ), .D(\R_DATA_TEMPR19[32] ), .Y(
        OR4_172_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C17 (.A_DOUT({
        nc8892, nc8893, nc8894, nc8895, nc8896, nc8897, nc8898, nc8899, 
        nc8900, nc8901, nc8902, nc8903, nc8904, nc8905, nc8906, nc8907, 
        nc8908, nc8909, \R_DATA_TEMPR14[35] , \R_DATA_TEMPR14[34] }), 
        .B_DOUT({nc8910, nc8911, nc8912, nc8913, nc8914, nc8915, 
        nc8916, nc8917, nc8918, nc8919, nc8920, nc8921, nc8922, nc8923, 
        nc8924, nc8925, nc8926, nc8927, nc8928, nc8929}), .DB_DETECT(
        \DB_DETECT[14][17] ), .SB_CORRECT(\SB_CORRECT[14][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C4 (.A_DOUT({nc8930, 
        nc8931, nc8932, nc8933, nc8934, nc8935, nc8936, nc8937, nc8938, 
        nc8939, nc8940, nc8941, nc8942, nc8943, nc8944, nc8945, nc8946, 
        nc8947, \R_DATA_TEMPR14[9] , \R_DATA_TEMPR14[8] }), .B_DOUT({
        nc8948, nc8949, nc8950, nc8951, nc8952, nc8953, nc8954, nc8955, 
        nc8956, nc8957, nc8958, nc8959, nc8960, nc8961, nc8962, nc8963, 
        nc8964, nc8965, nc8966, nc8967}), .DB_DETECT(
        \DB_DETECT[14][4] ), .SB_CORRECT(\SB_CORRECT[14][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C17 (.A_DOUT({
        nc8968, nc8969, nc8970, nc8971, nc8972, nc8973, nc8974, nc8975, 
        nc8976, nc8977, nc8978, nc8979, nc8980, nc8981, nc8982, nc8983, 
        nc8984, nc8985, \R_DATA_TEMPR30[35] , \R_DATA_TEMPR30[34] }), 
        .B_DOUT({nc8986, nc8987, nc8988, nc8989, nc8990, nc8991, 
        nc8992, nc8993, nc8994, nc8995, nc8996, nc8997, nc8998, nc8999, 
        nc9000, nc9001, nc9002, nc9003, nc9004, nc9005}), .DB_DETECT(
        \DB_DETECT[30][17] ), .SB_CORRECT(\SB_CORRECT[30][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_255 (.A(\R_DATA_TEMPR8[0] ), .B(\R_DATA_TEMPR9[0] ), .C(
        \R_DATA_TEMPR10[0] ), .D(\R_DATA_TEMPR11[0] ), .Y(OR4_255_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C8 (.A_DOUT({nc9006, 
        nc9007, nc9008, nc9009, nc9010, nc9011, nc9012, nc9013, nc9014, 
        nc9015, nc9016, nc9017, nc9018, nc9019, nc9020, nc9021, nc9022, 
        nc9023, \R_DATA_TEMPR17[17] , \R_DATA_TEMPR17[16] }), .B_DOUT({
        nc9024, nc9025, nc9026, nc9027, nc9028, nc9029, nc9030, nc9031, 
        nc9032, nc9033, nc9034, nc9035, nc9036, nc9037, nc9038, nc9039, 
        nc9040, nc9041, nc9042, nc9043}), .DB_DETECT(
        \DB_DETECT[17][8] ), .SB_CORRECT(\SB_CORRECT[17][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_190 (.A(\R_DATA_TEMPR8[8] ), .B(\R_DATA_TEMPR9[8] ), .C(
        \R_DATA_TEMPR10[8] ), .D(\R_DATA_TEMPR11[8] ), .Y(OR4_190_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C14 (.A_DOUT({
        nc9044, nc9045, nc9046, nc9047, nc9048, nc9049, nc9050, nc9051, 
        nc9052, nc9053, nc9054, nc9055, nc9056, nc9057, nc9058, nc9059, 
        nc9060, nc9061, \R_DATA_TEMPR12[29] , \R_DATA_TEMPR12[28] }), 
        .B_DOUT({nc9062, nc9063, nc9064, nc9065, nc9066, nc9067, 
        nc9068, nc9069, nc9070, nc9071, nc9072, nc9073, nc9074, nc9075, 
        nc9076, nc9077, nc9078, nc9079, nc9080, nc9081}), .DB_DETECT(
        \DB_DETECT[12][14] ), .SB_CORRECT(\SB_CORRECT[12][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C17 (.A_DOUT({
        nc9082, nc9083, nc9084, nc9085, nc9086, nc9087, nc9088, nc9089, 
        nc9090, nc9091, nc9092, nc9093, nc9094, nc9095, nc9096, nc9097, 
        nc9098, nc9099, \R_DATA_TEMPR15[35] , \R_DATA_TEMPR15[34] }), 
        .B_DOUT({nc9100, nc9101, nc9102, nc9103, nc9104, nc9105, 
        nc9106, nc9107, nc9108, nc9109, nc9110, nc9111, nc9112, nc9113, 
        nc9114, nc9115, nc9116, nc9117, nc9118, nc9119}), .DB_DETECT(
        \DB_DETECT[15][17] ), .SB_CORRECT(\SB_CORRECT[15][17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][17] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_26 (.A(OR4_189_Y), .B(OR2_28_Y), .C(\R_DATA_TEMPR22[19] ), 
        .D(\R_DATA_TEMPR23[19] ), .Y(OR4_26_Y));
    OR4 OR4_53 (.A(\R_DATA_TEMPR16[13] ), .B(\R_DATA_TEMPR17[13] ), .C(
        \R_DATA_TEMPR18[13] ), .D(\R_DATA_TEMPR19[13] ), .Y(OR4_53_Y));
    OR4 OR4_209 (.A(\R_DATA_TEMPR16[1] ), .B(\R_DATA_TEMPR17[1] ), .C(
        \R_DATA_TEMPR18[1] ), .D(\R_DATA_TEMPR19[1] ), .Y(OR4_209_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C14 (.A_DOUT({nc9120, 
        nc9121, nc9122, nc9123, nc9124, nc9125, nc9126, nc9127, nc9128, 
        nc9129, nc9130, nc9131, nc9132, nc9133, nc9134, nc9135, nc9136, 
        nc9137, \R_DATA_TEMPR5[29] , \R_DATA_TEMPR5[28] }), .B_DOUT({
        nc9138, nc9139, nc9140, nc9141, nc9142, nc9143, nc9144, nc9145, 
        nc9146, nc9147, nc9148, nc9149, nc9150, nc9151, nc9152, nc9153, 
        nc9154, nc9155, nc9156, nc9157}), .DB_DETECT(
        \DB_DETECT[5][14] ), .SB_CORRECT(\SB_CORRECT[5][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][14] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C4 (.A_DOUT({nc9158, 
        nc9159, nc9160, nc9161, nc9162, nc9163, nc9164, nc9165, nc9166, 
        nc9167, nc9168, nc9169, nc9170, nc9171, nc9172, nc9173, nc9174, 
        nc9175, \R_DATA_TEMPR26[9] , \R_DATA_TEMPR26[8] }), .B_DOUT({
        nc9176, nc9177, nc9178, nc9179, nc9180, nc9181, nc9182, nc9183, 
        nc9184, nc9185, nc9186, nc9187, nc9188, nc9189, nc9190, nc9191, 
        nc9192, nc9193, nc9194, nc9195}), .DB_DETECT(
        \DB_DETECT[26][4] ), .SB_CORRECT(\SB_CORRECT[26][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][4] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_279 (.A(\R_DATA_TEMPR28[9] ), .B(\R_DATA_TEMPR29[9] ), .C(
        \R_DATA_TEMPR30[9] ), .D(\R_DATA_TEMPR31[9] ), .Y(OR4_279_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C12 (.A_DOUT({
        nc9196, nc9197, nc9198, nc9199, nc9200, nc9201, nc9202, nc9203, 
        nc9204, nc9205, nc9206, nc9207, nc9208, nc9209, nc9210, nc9211, 
        nc9212, nc9213, \R_DATA_TEMPR26[25] , \R_DATA_TEMPR26[24] }), 
        .B_DOUT({nc9214, nc9215, nc9216, nc9217, nc9218, nc9219, 
        nc9220, nc9221, nc9222, nc9223, nc9224, nc9225, nc9226, nc9227, 
        nc9228, nc9229, nc9230, nc9231, nc9232, nc9233}), .DB_DETECT(
        \DB_DETECT[26][12] ), .SB_CORRECT(\SB_CORRECT[26][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C2 (.A_DOUT({nc9234, 
        nc9235, nc9236, nc9237, nc9238, nc9239, nc9240, nc9241, nc9242, 
        nc9243, nc9244, nc9245, nc9246, nc9247, nc9248, nc9249, nc9250, 
        nc9251, \R_DATA_TEMPR20[5] , \R_DATA_TEMPR20[4] }), .B_DOUT({
        nc9252, nc9253, nc9254, nc9255, nc9256, nc9257, nc9258, nc9259, 
        nc9260, nc9261, nc9262, nc9263, nc9264, nc9265, nc9266, nc9267, 
        nc9268, nc9269, nc9270, nc9271}), .DB_DETECT(
        \DB_DETECT[20][2] ), .SB_CORRECT(\SB_CORRECT[20][2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][2] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C10 (.A_DOUT({
        nc9272, nc9273, nc9274, nc9275, nc9276, nc9277, nc9278, nc9279, 
        nc9280, nc9281, nc9282, nc9283, nc9284, nc9285, nc9286, nc9287, 
        nc9288, nc9289, \R_DATA_TEMPR26[21] , \R_DATA_TEMPR26[20] }), 
        .B_DOUT({nc9290, nc9291, nc9292, nc9293, nc9294, nc9295, 
        nc9296, nc9297, nc9298, nc9299, nc9300, nc9301, nc9302, nc9303, 
        nc9304, nc9305, nc9306, nc9307, nc9308, nc9309}), .DB_DETECT(
        \DB_DETECT[26][10] ), .SB_CORRECT(\SB_CORRECT[26][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C18 (.A_DOUT({nc9310, 
        nc9311, nc9312, nc9313, nc9314, nc9315, nc9316, nc9317, nc9318, 
        nc9319, nc9320, nc9321, nc9322, nc9323, nc9324, nc9325, nc9326, 
        nc9327, \R_DATA_TEMPR2[37] , \R_DATA_TEMPR2[36] }), .B_DOUT({
        nc9328, nc9329, nc9330, nc9331, nc9332, nc9333, nc9334, nc9335, 
        nc9336, nc9337, nc9338, nc9339, nc9340, nc9341, nc9342, nc9343, 
        nc9344, nc9345, nc9346, nc9347}), .DB_DETECT(
        \DB_DETECT[2][18] ), .SB_CORRECT(\SB_CORRECT[2][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C19 (.A_DOUT({
        nc9348, nc9349, nc9350, nc9351, nc9352, nc9353, nc9354, nc9355, 
        nc9356, nc9357, nc9358, nc9359, nc9360, nc9361, nc9362, nc9363, 
        nc9364, nc9365, \R_DATA_TEMPR27[39] , \R_DATA_TEMPR27[38] }), 
        .B_DOUT({nc9366, nc9367, nc9368, nc9369, nc9370, nc9371, 
        nc9372, nc9373, nc9374, nc9375, nc9376, nc9377, nc9378, nc9379, 
        nc9380, nc9381, nc9382, nc9383, nc9384, nc9385}), .DB_DETECT(
        \DB_DETECT[27][19] ), .SB_CORRECT(\SB_CORRECT[27][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][19] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C6 (.A_DOUT({nc9386, 
        nc9387, nc9388, nc9389, nc9390, nc9391, nc9392, nc9393, nc9394, 
        nc9395, nc9396, nc9397, nc9398, nc9399, nc9400, nc9401, nc9402, 
        nc9403, \R_DATA_TEMPR14[13] , \R_DATA_TEMPR14[12] }), .B_DOUT({
        nc9404, nc9405, nc9406, nc9407, nc9408, nc9409, nc9410, nc9411, 
        nc9412, nc9413, nc9414, nc9415, nc9416, nc9417, nc9418, nc9419, 
        nc9420, nc9421, nc9422, nc9423}), .DB_DETECT(
        \DB_DETECT[14][6] ), .SB_CORRECT(\SB_CORRECT[14][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_89 (.A(OR4_110_Y), .B(OR4_221_Y), .C(OR4_316_Y), .D(
        OR4_123_Y), .Y(OR4_89_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C5 (.A_DOUT({nc9424, 
        nc9425, nc9426, nc9427, nc9428, nc9429, nc9430, nc9431, nc9432, 
        nc9433, nc9434, nc9435, nc9436, nc9437, nc9438, nc9439, nc9440, 
        nc9441, \R_DATA_TEMPR9[11] , \R_DATA_TEMPR9[10] }), .B_DOUT({
        nc9442, nc9443, nc9444, nc9445, nc9446, nc9447, nc9448, nc9449, 
        nc9450, nc9451, nc9452, nc9453, nc9454, nc9455, nc9456, nc9457, 
        nc9458, nc9459, nc9460, nc9461}), .DB_DETECT(\DB_DETECT[9][5] )
        , .SB_CORRECT(\SB_CORRECT[9][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_198 (.A(\R_DATA_TEMPR0[28] ), .B(\R_DATA_TEMPR1[28] ), .C(
        \R_DATA_TEMPR2[28] ), .D(\R_DATA_TEMPR3[28] ), .Y(OR4_198_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C10 (.A_DOUT({
        nc9462, nc9463, nc9464, nc9465, nc9466, nc9467, nc9468, nc9469, 
        nc9470, nc9471, nc9472, nc9473, nc9474, nc9475, nc9476, nc9477, 
        nc9478, nc9479, \R_DATA_TEMPR31[21] , \R_DATA_TEMPR31[20] }), 
        .B_DOUT({nc9480, nc9481, nc9482, nc9483, nc9484, nc9485, 
        nc9486, nc9487, nc9488, nc9489, nc9490, nc9491, nc9492, nc9493, 
        nc9494, nc9495, nc9496, nc9497, nc9498, nc9499}), .DB_DETECT(
        \DB_DETECT[31][10] ), .SB_CORRECT(\SB_CORRECT[31][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][10] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C5 (.A_DOUT({nc9500, 
        nc9501, nc9502, nc9503, nc9504, nc9505, nc9506, nc9507, nc9508, 
        nc9509, nc9510, nc9511, nc9512, nc9513, nc9514, nc9515, nc9516, 
        nc9517, \R_DATA_TEMPR19[11] , \R_DATA_TEMPR19[10] }), .B_DOUT({
        nc9518, nc9519, nc9520, nc9521, nc9522, nc9523, nc9524, nc9525, 
        nc9526, nc9527, nc9528, nc9529, nc9530, nc9531, nc9532, nc9533, 
        nc9534, nc9535, nc9536, nc9537}), .DB_DETECT(
        \DB_DETECT[19][5] ), .SB_CORRECT(\SB_CORRECT[19][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][5] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_258 (.A(\R_DATA_TEMPR8[13] ), .B(\R_DATA_TEMPR9[13] ), .C(
        \R_DATA_TEMPR10[13] ), .D(\R_DATA_TEMPR11[13] ), .Y(OR4_258_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_328_Y), .B(OR4_311_Y), .C(OR4_320_Y), 
        .D(OR4_202_Y), .Y(R_DATA[21]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C16 (.A_DOUT({nc9538, 
        nc9539, nc9540, nc9541, nc9542, nc9543, nc9544, nc9545, nc9546, 
        nc9547, nc9548, nc9549, nc9550, nc9551, nc9552, nc9553, nc9554, 
        nc9555, \R_DATA_TEMPR8[33] , \R_DATA_TEMPR8[32] }), .B_DOUT({
        nc9556, nc9557, nc9558, nc9559, nc9560, nc9561, nc9562, nc9563, 
        nc9564, nc9565, nc9566, nc9567, nc9568, nc9569, nc9570, nc9571, 
        nc9572, nc9573, nc9574, nc9575}), .DB_DETECT(
        \DB_DETECT[8][16] ), .SB_CORRECT(\SB_CORRECT[8][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C16 (.A_DOUT({
        nc9576, nc9577, nc9578, nc9579, nc9580, nc9581, nc9582, nc9583, 
        nc9584, nc9585, nc9586, nc9587, nc9588, nc9589, nc9590, nc9591, 
        nc9592, nc9593, \R_DATA_TEMPR16[33] , \R_DATA_TEMPR16[32] }), 
        .B_DOUT({nc9594, nc9595, nc9596, nc9597, nc9598, nc9599, 
        nc9600, nc9601, nc9602, nc9603, nc9604, nc9605, nc9606, nc9607, 
        nc9608, nc9609, nc9610, nc9611, nc9612, nc9613}), .DB_DETECT(
        \DB_DETECT[16][16] ), .SB_CORRECT(\SB_CORRECT[16][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][16] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_183 (.A(\R_DATA_TEMPR16[38] ), .B(\R_DATA_TEMPR17[38] ), 
        .C(\R_DATA_TEMPR18[38] ), .D(\R_DATA_TEMPR19[38] ), .Y(
        OR4_183_Y));
    OR4 OR4_332 (.A(\R_DATA_TEMPR8[32] ), .B(\R_DATA_TEMPR9[32] ), .C(
        \R_DATA_TEMPR10[32] ), .D(\R_DATA_TEMPR11[32] ), .Y(OR4_332_Y));
    OR4 OR4_247 (.A(\R_DATA_TEMPR8[12] ), .B(\R_DATA_TEMPR9[12] ), .C(
        \R_DATA_TEMPR10[12] ), .D(\R_DATA_TEMPR11[12] ), .Y(OR4_247_Y));
    OR4 OR4_13 (.A(OR4_67_Y), .B(OR2_4_Y), .C(\R_DATA_TEMPR22[10] ), 
        .D(\R_DATA_TEMPR23[10] ), .Y(OR4_13_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C6 (.A_DOUT({nc9614, 
        nc9615, nc9616, nc9617, nc9618, nc9619, nc9620, nc9621, nc9622, 
        nc9623, nc9624, nc9625, nc9626, nc9627, nc9628, nc9629, nc9630, 
        nc9631, \R_DATA_TEMPR22[13] , \R_DATA_TEMPR22[12] }), .B_DOUT({
        nc9632, nc9633, nc9634, nc9635, nc9636, nc9637, nc9638, nc9639, 
        nc9640, nc9641, nc9642, nc9643, nc9644, nc9645, nc9646, nc9647, 
        nc9648, nc9649, nc9650, nc9651}), .DB_DETECT(
        \DB_DETECT[22][6] ), .SB_CORRECT(\SB_CORRECT[22][6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][6] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C18 (.A_DOUT({nc9652, 
        nc9653, nc9654, nc9655, nc9656, nc9657, nc9658, nc9659, nc9660, 
        nc9661, nc9662, nc9663, nc9664, nc9665, nc9666, nc9667, nc9668, 
        nc9669, \R_DATA_TEMPR7[37] , \R_DATA_TEMPR7[36] }), .B_DOUT({
        nc9670, nc9671, nc9672, nc9673, nc9674, nc9675, nc9676, nc9677, 
        nc9678, nc9679, nc9680, nc9681, nc9682, nc9683, nc9684, nc9685, 
        nc9686, nc9687, nc9688, nc9689}), .DB_DETECT(
        \DB_DETECT[7][18] ), .SB_CORRECT(\SB_CORRECT[7][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_327 (.A(\R_DATA_TEMPR4[24] ), .B(\R_DATA_TEMPR5[24] ), .C(
        \R_DATA_TEMPR6[24] ), .D(\R_DATA_TEMPR7[24] ), .Y(OR4_327_Y));
    OR4 OR4_147 (.A(\R_DATA_TEMPR12[32] ), .B(\R_DATA_TEMPR13[32] ), 
        .C(\R_DATA_TEMPR14[32] ), .D(\R_DATA_TEMPR15[32] ), .Y(
        OR4_147_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C8 (.A_DOUT({nc9690, 
        nc9691, nc9692, nc9693, nc9694, nc9695, nc9696, nc9697, nc9698, 
        nc9699, nc9700, nc9701, nc9702, nc9703, nc9704, nc9705, nc9706, 
        nc9707, \R_DATA_TEMPR13[17] , \R_DATA_TEMPR13[16] }), .B_DOUT({
        nc9708, nc9709, nc9710, nc9711, nc9712, nc9713, nc9714, nc9715, 
        nc9716, nc9717, nc9718, nc9719, nc9720, nc9721, nc9722, nc9723, 
        nc9724, nc9725, nc9726, nc9727}), .DB_DETECT(
        \DB_DETECT[13][8] ), .SB_CORRECT(\SB_CORRECT[13][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][8] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_120 (.A(\R_DATA_TEMPR12[18] ), .B(\R_DATA_TEMPR13[18] ), 
        .C(\R_DATA_TEMPR14[18] ), .D(\R_DATA_TEMPR15[18] ), .Y(
        OR4_120_Y));
    OR4 OR4_51 (.A(OR4_157_Y), .B(OR4_288_Y), .C(OR4_252_Y), .D(
        OR4_112_Y), .Y(OR4_51_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C12 (.A_DOUT({
        nc9728, nc9729, nc9730, nc9731, nc9732, nc9733, nc9734, nc9735, 
        nc9736, nc9737, nc9738, nc9739, nc9740, nc9741, nc9742, nc9743, 
        nc9744, nc9745, \R_DATA_TEMPR10[25] , \R_DATA_TEMPR10[24] }), 
        .B_DOUT({nc9746, nc9747, nc9748, nc9749, nc9750, nc9751, 
        nc9752, nc9753, nc9754, nc9755, nc9756, nc9757, nc9758, nc9759, 
        nc9760, nc9761, nc9762, nc9763, nc9764, nc9765}), .DB_DETECT(
        \DB_DETECT[10][12] ), .SB_CORRECT(\SB_CORRECT[10][12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][12] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C11 (.A_DOUT({
        nc9766, nc9767, nc9768, nc9769, nc9770, nc9771, nc9772, nc9773, 
        nc9774, nc9775, nc9776, nc9777, nc9778, nc9779, nc9780, nc9781, 
        nc9782, nc9783, \R_DATA_TEMPR20[23] , \R_DATA_TEMPR20[22] }), 
        .B_DOUT({nc9784, nc9785, nc9786, nc9787, nc9788, nc9789, 
        nc9790, nc9791, nc9792, nc9793, nc9794, nc9795, nc9796, nc9797, 
        nc9798, nc9799, nc9800, nc9801, nc9802, nc9803}), .DB_DETECT(
        \DB_DETECT[20][11] ), .SB_CORRECT(\SB_CORRECT[20][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    INV \INVBLKY1[0]  (.A(R_ADDR[14]), .Y(\BLKY1[0] ));
    OR2 OR2_2 (.A(\R_DATA_TEMPR20[26] ), .B(\R_DATA_TEMPR21[26] ), .Y(
        OR2_2_Y));
    CFG2 #( .INIT(4'h8) )  CFG2_5 (.A(R_ADDR[16]), .B(R_ADDR[15]), .Y(
        CFG2_5_Y));
    OR4 \OR4_R_DATA[20]  (.A(OR4_262_Y), .B(OR4_351_Y), .C(OR4_141_Y), 
        .D(OR4_10_Y), .Y(R_DATA[20]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C6 (.A_DOUT({nc9804, 
        nc9805, nc9806, nc9807, nc9808, nc9809, nc9810, nc9811, nc9812, 
        nc9813, nc9814, nc9815, nc9816, nc9817, nc9818, nc9819, nc9820, 
        nc9821, \R_DATA_TEMPR0[13] , \R_DATA_TEMPR0[12] }), .B_DOUT({
        nc9822, nc9823, nc9824, nc9825, nc9826, nc9827, nc9828, nc9829, 
        nc9830, nc9831, nc9832, nc9833, nc9834, nc9835, nc9836, nc9837, 
        nc9838, nc9839, nc9840, nc9841}), .DB_DETECT(\DB_DETECT[0][6] )
        , .SB_CORRECT(\SB_CORRECT[0][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C11 (.A_DOUT({
        nc9842, nc9843, nc9844, nc9845, nc9846, nc9847, nc9848, nc9849, 
        nc9850, nc9851, nc9852, nc9853, nc9854, nc9855, nc9856, nc9857, 
        nc9858, nc9859, \R_DATA_TEMPR30[23] , \R_DATA_TEMPR30[22] }), 
        .B_DOUT({nc9860, nc9861, nc9862, nc9863, nc9864, nc9865, 
        nc9866, nc9867, nc9868, nc9869, nc9870, nc9871, nc9872, nc9873, 
        nc9874, nc9875, nc9876, nc9877, nc9878, nc9879}), .DB_DETECT(
        \DB_DETECT[30][11] ), .SB_CORRECT(\SB_CORRECT[30][11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][11] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C18 (.A_DOUT({
        nc9880, nc9881, nc9882, nc9883, nc9884, nc9885, nc9886, nc9887, 
        nc9888, nc9889, nc9890, nc9891, nc9892, nc9893, nc9894, nc9895, 
        nc9896, nc9897, \R_DATA_TEMPR27[37] , \R_DATA_TEMPR27[36] }), 
        .B_DOUT({nc9898, nc9899, nc9900, nc9901, nc9902, nc9903, 
        nc9904, nc9905, nc9906, nc9907, nc9908, nc9909, nc9910, nc9911, 
        nc9912, nc9913, nc9914, nc9915, nc9916, nc9917}), .DB_DETECT(
        \DB_DETECT[27][18] ), .SB_CORRECT(\SB_CORRECT[27][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_39 (.A(\R_DATA_TEMPR20[29] ), .B(\R_DATA_TEMPR21[29] ), .Y(
        OR2_39_Y));
    OR4 OR4_20 (.A(\R_DATA_TEMPR16[4] ), .B(\R_DATA_TEMPR17[4] ), .C(
        \R_DATA_TEMPR18[4] ), .D(\R_DATA_TEMPR19[4] ), .Y(OR4_20_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C3 (.A_DOUT({nc9918, 
        nc9919, nc9920, nc9921, nc9922, nc9923, nc9924, nc9925, nc9926, 
        nc9927, nc9928, nc9929, nc9930, nc9931, nc9932, nc9933, nc9934, 
        nc9935, \R_DATA_TEMPR5[7] , \R_DATA_TEMPR5[6] }), .B_DOUT({
        nc9936, nc9937, nc9938, nc9939, nc9940, nc9941, nc9942, nc9943, 
        nc9944, nc9945, nc9946, nc9947, nc9948, nc9949, nc9950, nc9951, 
        nc9952, nc9953, nc9954, nc9955}), .DB_DETECT(\DB_DETECT[5][3] )
        , .SB_CORRECT(\SB_CORRECT[5][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[26]  (.A(OR4_135_Y), .B(OR4_331_Y), .C(OR4_28_Y), 
        .D(OR4_48_Y), .Y(R_DATA[26]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C18 (.A_DOUT({
        nc9956, nc9957, nc9958, nc9959, nc9960, nc9961, nc9962, nc9963, 
        nc9964, nc9965, nc9966, nc9967, nc9968, nc9969, nc9970, nc9971, 
        nc9972, nc9973, \R_DATA_TEMPR30[37] , \R_DATA_TEMPR30[36] }), 
        .B_DOUT({nc9974, nc9975, nc9976, nc9977, nc9978, nc9979, 
        nc9980, nc9981, nc9982, nc9983, nc9984, nc9985, nc9986, nc9987, 
        nc9988, nc9989, nc9990, nc9991, nc9992, nc9993}), .DB_DETECT(
        \DB_DETECT[30][18] ), .SB_CORRECT(\SB_CORRECT[30][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][18] ), .A_ADDR({R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_244 (.A(OR4_195_Y), .B(OR2_24_Y), .C(\R_DATA_TEMPR22[17] ), 
        .D(\R_DATA_TEMPR23[17] ), .Y(OR4_244_Y));
    OR4 OR4_27 (.A(OR4_168_Y), .B(OR4_18_Y), .C(OR4_34_Y), .D(
        OR4_218_Y), .Y(OR4_27_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C13 (.A_DOUT({nc9994, 
        nc9995, nc9996, nc9997, nc9998, nc9999, nc10000, nc10001, 
        nc10002, nc10003, nc10004, nc10005, nc10006, nc10007, nc10008, 
        nc10009, nc10010, nc10011, \R_DATA_TEMPR4[27] , 
        \R_DATA_TEMPR4[26] }), .B_DOUT({nc10012, nc10013, nc10014, 
        nc10015, nc10016, nc10017, nc10018, nc10019, nc10020, nc10021, 
        nc10022, nc10023, nc10024, nc10025, nc10026, nc10027, nc10028, 
        nc10029, nc10030, nc10031}), .DB_DETECT(\DB_DETECT[4][13] ), 
        .SB_CORRECT(\SB_CORRECT[4][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_82 (.A(OR4_43_Y), .B(OR4_158_Y), .C(OR4_90_Y), .D(OR4_87_Y)
        , .Y(OR4_82_Y));
    OR4 OR4_230 (.A(\R_DATA_TEMPR24[25] ), .B(\R_DATA_TEMPR25[25] ), 
        .C(\R_DATA_TEMPR26[25] ), .D(\R_DATA_TEMPR27[25] ), .Y(
        OR4_230_Y));
    OR4 OR4_128 (.A(\R_DATA_TEMPR28[30] ), .B(\R_DATA_TEMPR29[30] ), 
        .C(\R_DATA_TEMPR30[30] ), .D(\R_DATA_TEMPR31[30] ), .Y(
        OR4_128_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1 (.A_DOUT({nc10032, 
        nc10033, nc10034, nc10035, nc10036, nc10037, nc10038, nc10039, 
        nc10040, nc10041, nc10042, nc10043, nc10044, nc10045, nc10046, 
        nc10047, nc10048, nc10049, \R_DATA_TEMPR3[3] , 
        \R_DATA_TEMPR3[2] }), .B_DOUT({nc10050, nc10051, nc10052, 
        nc10053, nc10054, nc10055, nc10056, nc10057, nc10058, nc10059, 
        nc10060, nc10061, nc10062, nc10063, nc10064, nc10065, nc10066, 
        nc10067, nc10068, nc10069}), .DB_DETECT(\DB_DETECT[3][1] ), 
        .SB_CORRECT(\SB_CORRECT[3][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C2 (.A_DOUT({
        nc10070, nc10071, nc10072, nc10073, nc10074, nc10075, nc10076, 
        nc10077, nc10078, nc10079, nc10080, nc10081, nc10082, nc10083, 
        nc10084, nc10085, nc10086, nc10087, \R_DATA_TEMPR16[5] , 
        \R_DATA_TEMPR16[4] }), .B_DOUT({nc10088, nc10089, nc10090, 
        nc10091, nc10092, nc10093, nc10094, nc10095, nc10096, nc10097, 
        nc10098, nc10099, nc10100, nc10101, nc10102, nc10103, nc10104, 
        nc10105, nc10106, nc10107}), .DB_DETECT(\DB_DETECT[16][2] ), 
        .SB_CORRECT(\SB_CORRECT[16][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C7 (.A_DOUT({
        nc10108, nc10109, nc10110, nc10111, nc10112, nc10113, nc10114, 
        nc10115, nc10116, nc10117, nc10118, nc10119, nc10120, nc10121, 
        nc10122, nc10123, nc10124, nc10125, \R_DATA_TEMPR16[15] , 
        \R_DATA_TEMPR16[14] }), .B_DOUT({nc10126, nc10127, nc10128, 
        nc10129, nc10130, nc10131, nc10132, nc10133, nc10134, nc10135, 
        nc10136, nc10137, nc10138, nc10139, nc10140, nc10141, nc10142, 
        nc10143, nc10144, nc10145}), .DB_DETECT(\DB_DETECT[16][7] ), 
        .SB_CORRECT(\SB_CORRECT[16][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C19 (.A_DOUT({
        nc10146, nc10147, nc10148, nc10149, nc10150, nc10151, nc10152, 
        nc10153, nc10154, nc10155, nc10156, nc10157, nc10158, nc10159, 
        nc10160, nc10161, nc10162, nc10163, \R_DATA_TEMPR22[39] , 
        \R_DATA_TEMPR22[38] }), .B_DOUT({nc10164, nc10165, nc10166, 
        nc10167, nc10168, nc10169, nc10170, nc10171, nc10172, nc10173, 
        nc10174, nc10175, nc10176, nc10177, nc10178, nc10179, nc10180, 
        nc10181, nc10182, nc10183}), .DB_DETECT(\DB_DETECT[22][19] ), 
        .SB_CORRECT(\SB_CORRECT[22][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C10 (.A_DOUT({
        nc10184, nc10185, nc10186, nc10187, nc10188, nc10189, nc10190, 
        nc10191, nc10192, nc10193, nc10194, nc10195, nc10196, nc10197, 
        nc10198, nc10199, nc10200, nc10201, \R_DATA_TEMPR11[21] , 
        \R_DATA_TEMPR11[20] }), .B_DOUT({nc10202, nc10203, nc10204, 
        nc10205, nc10206, nc10207, nc10208, nc10209, nc10210, nc10211, 
        nc10212, nc10213, nc10214, nc10215, nc10216, nc10217, nc10218, 
        nc10219, nc10220, nc10221}), .DB_DETECT(\DB_DETECT[11][10] ), 
        .SB_CORRECT(\SB_CORRECT[11][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_182 (.A(\R_DATA_TEMPR16[9] ), .B(\R_DATA_TEMPR17[9] ), .C(
        \R_DATA_TEMPR18[9] ), .D(\R_DATA_TEMPR19[9] ), .Y(OR4_182_Y));
    OR4 OR4_312 (.A(OR4_96_Y), .B(OR4_302_Y), .C(OR4_319_Y), .D(
        OR4_136_Y), .Y(OR4_312_Y));
    OR4 OR4_64 (.A(\R_DATA_TEMPR16[35] ), .B(\R_DATA_TEMPR17[35] ), .C(
        \R_DATA_TEMPR18[35] ), .D(\R_DATA_TEMPR19[35] ), .Y(OR4_64_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C13 (.A_DOUT({
        nc10222, nc10223, nc10224, nc10225, nc10226, nc10227, nc10228, 
        nc10229, nc10230, nc10231, nc10232, nc10233, nc10234, nc10235, 
        nc10236, nc10237, nc10238, nc10239, \R_DATA_TEMPR16[27] , 
        \R_DATA_TEMPR16[26] }), .B_DOUT({nc10240, nc10241, nc10242, 
        nc10243, nc10244, nc10245, nc10246, nc10247, nc10248, nc10249, 
        nc10250, nc10251, nc10252, nc10253, nc10254, nc10255, nc10256, 
        nc10257, nc10258, nc10259}), .DB_DETECT(\DB_DETECT[16][13] ), 
        .SB_CORRECT(\SB_CORRECT[16][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_11 (.A(\R_DATA_TEMPR24[6] ), .B(\R_DATA_TEMPR25[6] ), .C(
        \R_DATA_TEMPR26[6] ), .D(\R_DATA_TEMPR27[6] ), .Y(OR4_11_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C15 (.A_DOUT({
        nc10260, nc10261, nc10262, nc10263, nc10264, nc10265, nc10266, 
        nc10267, nc10268, nc10269, nc10270, nc10271, nc10272, nc10273, 
        nc10274, nc10275, nc10276, nc10277, \R_DATA_TEMPR11[31] , 
        \R_DATA_TEMPR11[30] }), .B_DOUT({nc10278, nc10279, nc10280, 
        nc10281, nc10282, nc10283, nc10284, nc10285, nc10286, nc10287, 
        nc10288, nc10289, nc10290, nc10291, nc10292, nc10293, nc10294, 
        nc10295, nc10296, nc10297}), .DB_DETECT(\DB_DETECT[11][15] ), 
        .SB_CORRECT(\SB_CORRECT[11][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C18 (.A_DOUT({
        nc10298, nc10299, nc10300, nc10301, nc10302, nc10303, nc10304, 
        nc10305, nc10306, nc10307, nc10308, nc10309, nc10310, nc10311, 
        nc10312, nc10313, nc10314, nc10315, \R_DATA_TEMPR5[37] , 
        \R_DATA_TEMPR5[36] }), .B_DOUT({nc10316, nc10317, nc10318, 
        nc10319, nc10320, nc10321, nc10322, nc10323, nc10324, nc10325, 
        nc10326, nc10327, nc10328, nc10329, nc10330, nc10331, nc10332, 
        nc10333, nc10334, nc10335}), .DB_DETECT(\DB_DETECT[5][18] ), 
        .SB_CORRECT(\SB_CORRECT[5][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C7 (.A_DOUT({
        nc10336, nc10337, nc10338, nc10339, nc10340, nc10341, nc10342, 
        nc10343, nc10344, nc10345, nc10346, nc10347, nc10348, nc10349, 
        nc10350, nc10351, nc10352, nc10353, \R_DATA_TEMPR12[15] , 
        \R_DATA_TEMPR12[14] }), .B_DOUT({nc10354, nc10355, nc10356, 
        nc10357, nc10358, nc10359, nc10360, nc10361, nc10362, nc10363, 
        nc10364, nc10365, nc10366, nc10367, nc10368, nc10369, nc10370, 
        nc10371, nc10372, nc10373}), .DB_DETECT(\DB_DETECT[12][7] ), 
        .SB_CORRECT(\SB_CORRECT[12][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C7 (.A_DOUT({nc10374, 
        nc10375, nc10376, nc10377, nc10378, nc10379, nc10380, nc10381, 
        nc10382, nc10383, nc10384, nc10385, nc10386, nc10387, nc10388, 
        nc10389, nc10390, nc10391, \R_DATA_TEMPR0[15] , 
        \R_DATA_TEMPR0[14] }), .B_DOUT({nc10392, nc10393, nc10394, 
        nc10395, nc10396, nc10397, nc10398, nc10399, nc10400, nc10401, 
        nc10402, nc10403, nc10404, nc10405, nc10406, nc10407, nc10408, 
        nc10409, nc10410, nc10411}), .DB_DETECT(\DB_DETECT[0][7] ), 
        .SB_CORRECT(\SB_CORRECT[0][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_345 (.A(OR4_42_Y), .B(OR4_257_Y), .C(OR4_332_Y), .D(
        OR4_147_Y), .Y(OR4_345_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C3 (.A_DOUT({nc10412, 
        nc10413, nc10414, nc10415, nc10416, nc10417, nc10418, nc10419, 
        nc10420, nc10421, nc10422, nc10423, nc10424, nc10425, nc10426, 
        nc10427, nc10428, nc10429, \R_DATA_TEMPR9[7] , 
        \R_DATA_TEMPR9[6] }), .B_DOUT({nc10430, nc10431, nc10432, 
        nc10433, nc10434, nc10435, nc10436, nc10437, nc10438, nc10439, 
        nc10440, nc10441, nc10442, nc10443, nc10444, nc10445, nc10446, 
        nc10447, nc10448, nc10449}), .DB_DETECT(\DB_DETECT[9][3] ), 
        .SB_CORRECT(\SB_CORRECT[9][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_236 (.A(\R_DATA_TEMPR24[1] ), .B(\R_DATA_TEMPR25[1] ), .C(
        \R_DATA_TEMPR26[1] ), .D(\R_DATA_TEMPR27[1] ), .Y(OR4_236_Y));
    OR2 OR2_7 (.A(\R_DATA_TEMPR20[15] ), .B(\R_DATA_TEMPR21[15] ), .Y(
        OR2_7_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C12 (.A_DOUT({
        nc10450, nc10451, nc10452, nc10453, nc10454, nc10455, nc10456, 
        nc10457, nc10458, nc10459, nc10460, nc10461, nc10462, nc10463, 
        nc10464, nc10465, nc10466, nc10467, \R_DATA_TEMPR14[25] , 
        \R_DATA_TEMPR14[24] }), .B_DOUT({nc10468, nc10469, nc10470, 
        nc10471, nc10472, nc10473, nc10474, nc10475, nc10476, nc10477, 
        nc10478, nc10479, nc10480, nc10481, nc10482, nc10483, nc10484, 
        nc10485, nc10486, nc10487}), .DB_DETECT(\DB_DETECT[14][12] ), 
        .SB_CORRECT(\SB_CORRECT[14][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C11 (.A_DOUT({
        nc10488, nc10489, nc10490, nc10491, nc10492, nc10493, nc10494, 
        nc10495, nc10496, nc10497, nc10498, nc10499, nc10500, nc10501, 
        nc10502, nc10503, nc10504, nc10505, \R_DATA_TEMPR24[23] , 
        \R_DATA_TEMPR24[22] }), .B_DOUT({nc10506, nc10507, nc10508, 
        nc10509, nc10510, nc10511, nc10512, nc10513, nc10514, nc10515, 
        nc10516, nc10517, nc10518, nc10519, nc10520, nc10521, nc10522, 
        nc10523, nc10524, nc10525}), .DB_DETECT(\DB_DETECT[24][11] ), 
        .SB_CORRECT(\SB_CORRECT[24][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C17 (.A_DOUT({
        nc10526, nc10527, nc10528, nc10529, nc10530, nc10531, nc10532, 
        nc10533, nc10534, nc10535, nc10536, nc10537, nc10538, nc10539, 
        nc10540, nc10541, nc10542, nc10543, \R_DATA_TEMPR3[35] , 
        \R_DATA_TEMPR3[34] }), .B_DOUT({nc10544, nc10545, nc10546, 
        nc10547, nc10548, nc10549, nc10550, nc10551, nc10552, nc10553, 
        nc10554, nc10555, nc10556, nc10557, nc10558, nc10559, nc10560, 
        nc10561, nc10562, nc10563}), .DB_DETECT(\DB_DETECT[3][17] ), 
        .SB_CORRECT(\SB_CORRECT[3][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_73 (.A(\R_DATA_TEMPR12[10] ), .B(\R_DATA_TEMPR13[10] ), .C(
        \R_DATA_TEMPR14[10] ), .D(\R_DATA_TEMPR15[10] ), .Y(OR4_73_Y));
    OR4 OR4_195 (.A(\R_DATA_TEMPR16[17] ), .B(\R_DATA_TEMPR17[17] ), 
        .C(\R_DATA_TEMPR18[17] ), .D(\R_DATA_TEMPR19[17] ), .Y(
        OR4_195_Y));
    OR4 OR4_252 (.A(\R_DATA_TEMPR8[5] ), .B(\R_DATA_TEMPR9[5] ), .C(
        \R_DATA_TEMPR10[5] ), .D(\R_DATA_TEMPR11[5] ), .Y(OR4_252_Y));
    OR4 OR4_289 (.A(\R_DATA_TEMPR12[26] ), .B(\R_DATA_TEMPR13[26] ), 
        .C(\R_DATA_TEMPR14[26] ), .D(\R_DATA_TEMPR15[26] ), .Y(
        OR4_289_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C17 (.A_DOUT({
        nc10564, nc10565, nc10566, nc10567, nc10568, nc10569, nc10570, 
        nc10571, nc10572, nc10573, nc10574, nc10575, nc10576, nc10577, 
        nc10578, nc10579, nc10580, nc10581, \R_DATA_TEMPR26[35] , 
        \R_DATA_TEMPR26[34] }), .B_DOUT({nc10582, nc10583, nc10584, 
        nc10585, nc10586, nc10587, nc10588, nc10589, nc10590, nc10591, 
        nc10592, nc10593, nc10594, nc10595, nc10596, nc10597, nc10598, 
        nc10599, nc10600, nc10601}), .DB_DETECT(\DB_DETECT[26][17] ), 
        .SB_CORRECT(\SB_CORRECT[26][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_32 (.A(\R_DATA_TEMPR20[39] ), .B(\R_DATA_TEMPR21[39] ), .Y(
        OR2_32_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C12 (.A_DOUT({
        nc10602, nc10603, nc10604, nc10605, nc10606, nc10607, nc10608, 
        nc10609, nc10610, nc10611, nc10612, nc10613, nc10614, nc10615, 
        nc10616, nc10617, nc10618, nc10619, \R_DATA_TEMPR27[25] , 
        \R_DATA_TEMPR27[24] }), .B_DOUT({nc10620, nc10621, nc10622, 
        nc10623, nc10624, nc10625, nc10626, nc10627, nc10628, nc10629, 
        nc10630, nc10631, nc10632, nc10633, nc10634, nc10635, nc10636, 
        nc10637, nc10638, nc10639}), .DB_DETECT(\DB_DETECT[27][12] ), 
        .SB_CORRECT(\SB_CORRECT[27][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C11 (.A_DOUT({
        nc10640, nc10641, nc10642, nc10643, nc10644, nc10645, nc10646, 
        nc10647, nc10648, nc10649, nc10650, nc10651, nc10652, nc10653, 
        nc10654, nc10655, nc10656, nc10657, \R_DATA_TEMPR25[23] , 
        \R_DATA_TEMPR25[22] }), .B_DOUT({nc10658, nc10659, nc10660, 
        nc10661, nc10662, nc10663, nc10664, nc10665, nc10666, nc10667, 
        nc10668, nc10669, nc10670, nc10671, nc10672, nc10673, nc10674, 
        nc10675, nc10676, nc10677}), .DB_DETECT(\DB_DETECT[25][11] ), 
        .SB_CORRECT(\SB_CORRECT[25][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C12 (.A_DOUT({
        nc10678, nc10679, nc10680, nc10681, nc10682, nc10683, nc10684, 
        nc10685, nc10686, nc10687, nc10688, nc10689, nc10690, nc10691, 
        nc10692, nc10693, nc10694, nc10695, \R_DATA_TEMPR15[25] , 
        \R_DATA_TEMPR15[24] }), .B_DOUT({nc10696, nc10697, nc10698, 
        nc10699, nc10700, nc10701, nc10702, nc10703, nc10704, nc10705, 
        nc10706, nc10707, nc10708, nc10709, nc10710, nc10711, nc10712, 
        nc10713, nc10714, nc10715}), .DB_DETECT(\DB_DETECT[15][12] ), 
        .SB_CORRECT(\SB_CORRECT[15][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C10 (.A_DOUT({
        nc10716, nc10717, nc10718, nc10719, nc10720, nc10721, nc10722, 
        nc10723, nc10724, nc10725, nc10726, nc10727, nc10728, nc10729, 
        nc10730, nc10731, nc10732, nc10733, \R_DATA_TEMPR27[21] , 
        \R_DATA_TEMPR27[20] }), .B_DOUT({nc10734, nc10735, nc10736, 
        nc10737, nc10738, nc10739, nc10740, nc10741, nc10742, nc10743, 
        nc10744, nc10745, nc10746, nc10747, nc10748, nc10749, nc10750, 
        nc10751, nc10752, nc10753}), .DB_DETECT(\DB_DETECT[27][10] ), 
        .SB_CORRECT(\SB_CORRECT[27][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_1 (.A(\R_DATA_TEMPR20[33] ), .B(\R_DATA_TEMPR21[33] ), .Y(
        OR2_1_Y));
    OR4 OR4_210 (.A(OR4_309_Y), .B(OR2_12_Y), .C(\R_DATA_TEMPR22[14] ), 
        .D(\R_DATA_TEMPR23[14] ), .Y(OR4_210_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C18 (.A_DOUT({
        nc10754, nc10755, nc10756, nc10757, nc10758, nc10759, nc10760, 
        nc10761, nc10762, nc10763, nc10764, nc10765, nc10766, nc10767, 
        nc10768, nc10769, nc10770, nc10771, \R_DATA_TEMPR22[37] , 
        \R_DATA_TEMPR22[36] }), .B_DOUT({nc10772, nc10773, nc10774, 
        nc10775, nc10776, nc10777, nc10778, nc10779, nc10780, nc10781, 
        nc10782, nc10783, nc10784, nc10785, nc10786, nc10787, nc10788, 
        nc10789, nc10790, nc10791}), .DB_DETECT(\DB_DETECT[22][18] ), 
        .SB_CORRECT(\SB_CORRECT[22][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C15 (.A_DOUT({
        nc10792, nc10793, nc10794, nc10795, nc10796, nc10797, nc10798, 
        nc10799, nc10800, nc10801, nc10802, nc10803, nc10804, nc10805, 
        nc10806, nc10807, nc10808, nc10809, \R_DATA_TEMPR9[31] , 
        \R_DATA_TEMPR9[30] }), .B_DOUT({nc10810, nc10811, nc10812, 
        nc10813, nc10814, nc10815, nc10816, nc10817, nc10818, nc10819, 
        nc10820, nc10821, nc10822, nc10823, nc10824, nc10825, nc10826, 
        nc10827, nc10828, nc10829}), .DB_DETECT(\DB_DETECT[9][15] ), 
        .SB_CORRECT(\SB_CORRECT[9][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C3 (.A_DOUT({
        nc10830, nc10831, nc10832, nc10833, nc10834, nc10835, nc10836, 
        nc10837, nc10838, nc10839, nc10840, nc10841, nc10842, nc10843, 
        nc10844, nc10845, nc10846, nc10847, \R_DATA_TEMPR14[7] , 
        \R_DATA_TEMPR14[6] }), .B_DOUT({nc10848, nc10849, nc10850, 
        nc10851, nc10852, nc10853, nc10854, nc10855, nc10856, nc10857, 
        nc10858, nc10859, nc10860, nc10861, nc10862, nc10863, nc10864, 
        nc10865, nc10866, nc10867}), .DB_DETECT(\DB_DETECT[14][3] ), 
        .SB_CORRECT(\SB_CORRECT[14][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_350 (.A(\R_DATA_TEMPR0[7] ), .B(\R_DATA_TEMPR1[7] ), .C(
        \R_DATA_TEMPR2[7] ), .D(\R_DATA_TEMPR3[7] ), .Y(OR4_350_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C9 (.A_DOUT({
        nc10868, nc10869, nc10870, nc10871, nc10872, nc10873, nc10874, 
        nc10875, nc10876, nc10877, nc10878, nc10879, nc10880, nc10881, 
        nc10882, nc10883, nc10884, nc10885, \R_DATA_TEMPR10[19] , 
        \R_DATA_TEMPR10[18] }), .B_DOUT({nc10886, nc10887, nc10888, 
        nc10889, nc10890, nc10891, nc10892, nc10893, nc10894, nc10895, 
        nc10896, nc10897, nc10898, nc10899, nc10900, nc10901, nc10902, 
        nc10903, nc10904, nc10905}), .DB_DETECT(\DB_DETECT[10][9] ), 
        .SB_CORRECT(\SB_CORRECT[10][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_295 (.A(OR4_108_Y), .B(OR2_13_Y), .C(\R_DATA_TEMPR22[18] ), 
        .D(\R_DATA_TEMPR23[18] ), .Y(OR4_295_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C5 (.A_DOUT({
        nc10906, nc10907, nc10908, nc10909, nc10910, nc10911, nc10912, 
        nc10913, nc10914, nc10915, nc10916, nc10917, nc10918, nc10919, 
        nc10920, nc10921, nc10922, nc10923, \R_DATA_TEMPR30[11] , 
        \R_DATA_TEMPR30[10] }), .B_DOUT({nc10924, nc10925, nc10926, 
        nc10927, nc10928, nc10929, nc10930, nc10931, nc10932, nc10933, 
        nc10934, nc10935, nc10936, nc10937, nc10938, nc10939, nc10940, 
        nc10941, nc10942, nc10943}), .DB_DETECT(\DB_DETECT[30][5] ), 
        .SB_CORRECT(\SB_CORRECT[30][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C16 (.A_DOUT({
        nc10944, nc10945, nc10946, nc10947, nc10948, nc10949, nc10950, 
        nc10951, nc10952, nc10953, nc10954, nc10955, nc10956, nc10957, 
        nc10958, nc10959, nc10960, nc10961, \R_DATA_TEMPR17[33] , 
        \R_DATA_TEMPR17[32] }), .B_DOUT({nc10962, nc10963, nc10964, 
        nc10965, nc10966, nc10967, nc10968, nc10969, nc10970, nc10971, 
        nc10972, nc10973, nc10974, nc10975, nc10976, nc10977, nc10978, 
        nc10979, nc10980, nc10981}), .DB_DETECT(\DB_DETECT[17][16] ), 
        .SB_CORRECT(\SB_CORRECT[17][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C14 (.A_DOUT({
        nc10982, nc10983, nc10984, nc10985, nc10986, nc10987, nc10988, 
        nc10989, nc10990, nc10991, nc10992, nc10993, nc10994, nc10995, 
        nc10996, nc10997, nc10998, nc10999, \R_DATA_TEMPR1[29] , 
        \R_DATA_TEMPR1[28] }), .B_DOUT({nc11000, nc11001, nc11002, 
        nc11003, nc11004, nc11005, nc11006, nc11007, nc11008, nc11009, 
        nc11010, nc11011, nc11012, nc11013, nc11014, nc11015, nc11016, 
        nc11017, nc11018, nc11019}), .DB_DETECT(\DB_DETECT[1][14] ), 
        .SB_CORRECT(\SB_CORRECT[1][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C12 (.A_DOUT({
        nc11020, nc11021, nc11022, nc11023, nc11024, nc11025, nc11026, 
        nc11027, nc11028, nc11029, nc11030, nc11031, nc11032, nc11033, 
        nc11034, nc11035, nc11036, nc11037, \R_DATA_TEMPR6[25] , 
        \R_DATA_TEMPR6[24] }), .B_DOUT({nc11038, nc11039, nc11040, 
        nc11041, nc11042, nc11043, nc11044, nc11045, nc11046, nc11047, 
        nc11048, nc11049, nc11050, nc11051, nc11052, nc11053, nc11054, 
        nc11055, nc11056, nc11057}), .DB_DETECT(\DB_DETECT[6][12] ), 
        .SB_CORRECT(\SB_CORRECT[6][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C14 (.A_DOUT({
        nc11058, nc11059, nc11060, nc11061, nc11062, nc11063, nc11064, 
        nc11065, nc11066, nc11067, nc11068, nc11069, nc11070, nc11071, 
        nc11072, nc11073, nc11074, nc11075, \R_DATA_TEMPR19[29] , 
        \R_DATA_TEMPR19[28] }), .B_DOUT({nc11076, nc11077, nc11078, 
        nc11079, nc11080, nc11081, nc11082, nc11083, nc11084, nc11085, 
        nc11086, nc11087, nc11088, nc11089, nc11090, nc11091, nc11092, 
        nc11093, nc11094, nc11095}), .DB_DETECT(\DB_DETECT[19][14] ), 
        .SB_CORRECT(\SB_CORRECT[19][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_35 (.A(\R_DATA_TEMPR0[4] ), .B(\R_DATA_TEMPR1[4] ), .C(
        \R_DATA_TEMPR2[4] ), .D(\R_DATA_TEMPR3[4] ), .Y(OR4_35_Y));
    OR4 OR4_216 (.A(\R_DATA_TEMPR8[22] ), .B(\R_DATA_TEMPR9[22] ), .C(
        \R_DATA_TEMPR10[22] ), .D(\R_DATA_TEMPR11[22] ), .Y(OR4_216_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C6 (.A_DOUT({
        nc11096, nc11097, nc11098, nc11099, nc11100, nc11101, nc11102, 
        nc11103, nc11104, nc11105, nc11106, nc11107, nc11108, nc11109, 
        nc11110, nc11111, nc11112, nc11113, \R_DATA_TEMPR10[13] , 
        \R_DATA_TEMPR10[12] }), .B_DOUT({nc11114, nc11115, nc11116, 
        nc11117, nc11118, nc11119, nc11120, nc11121, nc11122, nc11123, 
        nc11124, nc11125, nc11126, nc11127, nc11128, nc11129, nc11130, 
        nc11131, nc11132, nc11133}), .DB_DETECT(\DB_DETECT[10][6] ), 
        .SB_CORRECT(\SB_CORRECT[10][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C14 (.A_DOUT({
        nc11134, nc11135, nc11136, nc11137, nc11138, nc11139, nc11140, 
        nc11141, nc11142, nc11143, nc11144, nc11145, nc11146, nc11147, 
        nc11148, nc11149, nc11150, nc11151, \R_DATA_TEMPR26[29] , 
        \R_DATA_TEMPR26[28] }), .B_DOUT({nc11152, nc11153, nc11154, 
        nc11155, nc11156, nc11157, nc11158, nc11159, nc11160, nc11161, 
        nc11162, nc11163, nc11164, nc11165, nc11166, nc11167, nc11168, 
        nc11169, nc11170, nc11171}), .DB_DETECT(\DB_DETECT[26][14] ), 
        .SB_CORRECT(\SB_CORRECT[26][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_71 (.A(\R_DATA_TEMPR12[8] ), .B(\R_DATA_TEMPR13[8] ), .C(
        \R_DATA_TEMPR14[8] ), .D(\R_DATA_TEMPR15[8] ), .Y(OR4_71_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0 (.A_DOUT({
        nc11172, nc11173, nc11174, nc11175, nc11176, nc11177, nc11178, 
        nc11179, nc11180, nc11181, nc11182, nc11183, nc11184, nc11185, 
        nc11186, nc11187, nc11188, nc11189, \R_DATA_TEMPR31[1] , 
        \R_DATA_TEMPR31[0] }), .B_DOUT({nc11190, nc11191, nc11192, 
        nc11193, nc11194, nc11195, nc11196, nc11197, nc11198, nc11199, 
        nc11200, nc11201, nc11202, nc11203, nc11204, nc11205, nc11206, 
        nc11207, nc11208, nc11209}), .DB_DETECT(\DB_DETECT[31][0] ), 
        .SB_CORRECT(\SB_CORRECT[31][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_125 (.A(\R_DATA_TEMPR8[34] ), .B(\R_DATA_TEMPR9[34] ), .C(
        \R_DATA_TEMPR10[34] ), .D(\R_DATA_TEMPR11[34] ), .Y(OR4_125_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C9 (.A_DOUT({
        nc11210, nc11211, nc11212, nc11213, nc11214, nc11215, nc11216, 
        nc11217, nc11218, nc11219, nc11220, nc11221, nc11222, nc11223, 
        nc11224, nc11225, nc11226, nc11227, \R_DATA_TEMPR24[19] , 
        \R_DATA_TEMPR24[18] }), .B_DOUT({nc11228, nc11229, nc11230, 
        nc11231, nc11232, nc11233, nc11234, nc11235, nc11236, nc11237, 
        nc11238, nc11239, nc11240, nc11241, nc11242, nc11243, nc11244, 
        nc11245, nc11246, nc11247}), .DB_DETECT(\DB_DETECT[24][9] ), 
        .SB_CORRECT(\SB_CORRECT[24][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_298 (.A(\R_DATA_TEMPR28[5] ), .B(\R_DATA_TEMPR29[5] ), .C(
        \R_DATA_TEMPR30[5] ), .D(\R_DATA_TEMPR31[5] ), .Y(OR4_298_Y));
    OR4 \OR4_R_DATA[27]  (.A(OR4_40_Y), .B(OR4_211_Y), .C(OR4_306_Y), 
        .D(OR4_347_Y), .Y(R_DATA[27]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C19 (.A_DOUT({
        nc11248, nc11249, nc11250, nc11251, nc11252, nc11253, nc11254, 
        nc11255, nc11256, nc11257, nc11258, nc11259, nc11260, nc11261, 
        nc11262, nc11263, nc11264, nc11265, \R_DATA_TEMPR30[39] , 
        \R_DATA_TEMPR30[38] }), .B_DOUT({nc11266, nc11267, nc11268, 
        nc11269, nc11270, nc11271, nc11272, nc11273, nc11274, nc11275, 
        nc11276, nc11277, nc11278, nc11279, nc11280, nc11281, nc11282, 
        nc11283, nc11284, nc11285}), .DB_DETECT(\DB_DETECT[30][19] ), 
        .SB_CORRECT(\SB_CORRECT[30][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C11 (.A_DOUT({
        nc11286, nc11287, nc11288, nc11289, nc11290, nc11291, nc11292, 
        nc11293, nc11294, nc11295, nc11296, nc11297, nc11298, nc11299, 
        nc11300, nc11301, nc11302, nc11303, \R_DATA_TEMPR2[23] , 
        \R_DATA_TEMPR2[22] }), .B_DOUT({nc11304, nc11305, nc11306, 
        nc11307, nc11308, nc11309, nc11310, nc11311, nc11312, nc11313, 
        nc11314, nc11315, nc11316, nc11317, nc11318, nc11319, nc11320, 
        nc11321, nc11322, nc11323}), .DB_DETECT(\DB_DETECT[2][11] ), 
        .SB_CORRECT(\SB_CORRECT[2][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_28 (.A(\R_DATA_TEMPR24[26] ), .B(\R_DATA_TEMPR25[26] ), .C(
        \R_DATA_TEMPR26[26] ), .D(\R_DATA_TEMPR27[26] ), .Y(OR4_28_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C12 (.A_DOUT({
        nc11324, nc11325, nc11326, nc11327, nc11328, nc11329, nc11330, 
        nc11331, nc11332, nc11333, nc11334, nc11335, nc11336, nc11337, 
        nc11338, nc11339, nc11340, nc11341, \R_DATA_TEMPR22[25] , 
        \R_DATA_TEMPR22[24] }), .B_DOUT({nc11342, nc11343, nc11344, 
        nc11345, nc11346, nc11347, nc11348, nc11349, nc11350, nc11351, 
        nc11352, nc11353, nc11354, nc11355, nc11356, nc11357, nc11358, 
        nc11359, nc11360, nc11361}), .DB_DETECT(\DB_DETECT[22][12] ), 
        .SB_CORRECT(\SB_CORRECT[22][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C7 (.A_DOUT({
        nc11362, nc11363, nc11364, nc11365, nc11366, nc11367, nc11368, 
        nc11369, nc11370, nc11371, nc11372, nc11373, nc11374, nc11375, 
        nc11376, nc11377, nc11378, nc11379, \R_DATA_TEMPR17[15] , 
        \R_DATA_TEMPR17[14] }), .B_DOUT({nc11380, nc11381, nc11382, 
        nc11383, nc11384, nc11385, nc11386, nc11387, nc11388, nc11389, 
        nc11390, nc11391, nc11392, nc11393, nc11394, nc11395, nc11396, 
        nc11397, nc11398, nc11399}), .DB_DETECT(\DB_DETECT[17][7] ), 
        .SB_CORRECT(\SB_CORRECT[17][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[6]  (.A(CFG2_1_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[6] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C10 (.A_DOUT({
        nc11400, nc11401, nc11402, nc11403, nc11404, nc11405, nc11406, 
        nc11407, nc11408, nc11409, nc11410, nc11411, nc11412, nc11413, 
        nc11414, nc11415, nc11416, nc11417, \R_DATA_TEMPR22[21] , 
        \R_DATA_TEMPR22[20] }), .B_DOUT({nc11418, nc11419, nc11420, 
        nc11421, nc11422, nc11423, nc11424, nc11425, nc11426, nc11427, 
        nc11428, nc11429, nc11430, nc11431, nc11432, nc11433, nc11434, 
        nc11435, nc11436, nc11437}), .DB_DETECT(\DB_DETECT[22][10] ), 
        .SB_CORRECT(\SB_CORRECT[22][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_164 (.A(\R_DATA_TEMPR16[36] ), .B(\R_DATA_TEMPR17[36] ), 
        .C(\R_DATA_TEMPR18[36] ), .D(\R_DATA_TEMPR19[36] ), .Y(
        OR4_164_Y));
    OR4 OR4_225 (.A(OR4_296_Y), .B(OR4_140_Y), .C(OR4_216_Y), .D(
        OR4_36_Y), .Y(OR4_225_Y));
    CFG2 #( .INIT(4'h4) )  CFG2_2 (.A(W_ADDR[16]), .B(W_ADDR[15]), .Y(
        CFG2_2_Y));
    OR4 OR4_347 (.A(\R_DATA_TEMPR28[27] ), .B(\R_DATA_TEMPR29[27] ), 
        .C(\R_DATA_TEMPR30[27] ), .D(\R_DATA_TEMPR31[27] ), .Y(
        OR4_347_Y));
    OR4 OR4_140 (.A(\R_DATA_TEMPR4[22] ), .B(\R_DATA_TEMPR5[22] ), .C(
        \R_DATA_TEMPR6[22] ), .D(\R_DATA_TEMPR7[22] ), .Y(OR4_140_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C3 (.A_DOUT({
        nc11438, nc11439, nc11440, nc11441, nc11442, nc11443, nc11444, 
        nc11445, nc11446, nc11447, nc11448, nc11449, nc11450, nc11451, 
        nc11452, nc11453, nc11454, nc11455, \R_DATA_TEMPR11[7] , 
        \R_DATA_TEMPR11[6] }), .B_DOUT({nc11456, nc11457, nc11458, 
        nc11459, nc11460, nc11461, nc11462, nc11463, nc11464, nc11465, 
        nc11466, nc11467, nc11468, nc11469, nc11470, nc11471, nc11472, 
        nc11473, nc11474, nc11475}), .DB_DETECT(\DB_DETECT[11][3] ), 
        .SB_CORRECT(\SB_CORRECT[11][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C13 (.A_DOUT({
        nc11476, nc11477, nc11478, nc11479, nc11480, nc11481, nc11482, 
        nc11483, nc11484, nc11485, nc11486, nc11487, nc11488, nc11489, 
        nc11490, nc11491, nc11492, nc11493, \R_DATA_TEMPR17[27] , 
        \R_DATA_TEMPR17[26] }), .B_DOUT({nc11494, nc11495, nc11496, 
        nc11497, nc11498, nc11499, nc11500, nc11501, nc11502, nc11503, 
        nc11504, nc11505, nc11506, nc11507, nc11508, nc11509, nc11510, 
        nc11511, nc11512, nc11513}), .DB_DETECT(\DB_DETECT[17][13] ), 
        .SB_CORRECT(\SB_CORRECT[17][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C14 (.A_DOUT({
        nc11514, nc11515, nc11516, nc11517, nc11518, nc11519, nc11520, 
        nc11521, nc11522, nc11523, nc11524, nc11525, nc11526, nc11527, 
        nc11528, nc11529, nc11530, nc11531, \R_DATA_TEMPR8[29] , 
        \R_DATA_TEMPR8[28] }), .B_DOUT({nc11532, nc11533, nc11534, 
        nc11535, nc11536, nc11537, nc11538, nc11539, nc11540, nc11541, 
        nc11542, nc11543, nc11544, nc11545, nc11546, nc11547, nc11548, 
        nc11549, nc11550, nc11551}), .DB_DETECT(\DB_DETECT[8][14] ), 
        .SB_CORRECT(\SB_CORRECT[8][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_306 (.A(\R_DATA_TEMPR24[27] ), .B(\R_DATA_TEMPR25[27] ), 
        .C(\R_DATA_TEMPR26[27] ), .D(\R_DATA_TEMPR27[27] ), .Y(
        OR4_306_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C14 (.A_DOUT({
        nc11552, nc11553, nc11554, nc11555, nc11556, nc11557, nc11558, 
        nc11559, nc11560, nc11561, nc11562, nc11563, nc11564, nc11565, 
        nc11566, nc11567, nc11568, nc11569, \R_DATA_TEMPR31[29] , 
        \R_DATA_TEMPR31[28] }), .B_DOUT({nc11570, nc11571, nc11572, 
        nc11573, nc11574, nc11575, nc11576, nc11577, nc11578, nc11579, 
        nc11580, nc11581, nc11582, nc11583, nc11584, nc11585, nc11586, 
        nc11587, nc11588, nc11589}), .DB_DETECT(\DB_DETECT[31][14] ), 
        .SB_CORRECT(\SB_CORRECT[31][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C16 (.A_DOUT({
        nc11590, nc11591, nc11592, nc11593, nc11594, nc11595, nc11596, 
        nc11597, nc11598, nc11599, nc11600, nc11601, nc11602, nc11603, 
        nc11604, nc11605, nc11606, nc11607, \R_DATA_TEMPR12[33] , 
        \R_DATA_TEMPR12[32] }), .B_DOUT({nc11608, nc11609, nc11610, 
        nc11611, nc11612, nc11613, nc11614, nc11615, nc11616, nc11617, 
        nc11618, nc11619, nc11620, nc11621, nc11622, nc11623, nc11624, 
        nc11625, nc11626, nc11627}), .DB_DETECT(\DB_DETECT[12][16] ), 
        .SB_CORRECT(\SB_CORRECT[12][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h1) )  CFG2_3 (.A(R_ADDR[16]), .B(R_ADDR[15]), .Y(
        CFG2_3_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C11 (.A_DOUT({
        nc11628, nc11629, nc11630, nc11631, nc11632, nc11633, nc11634, 
        nc11635, nc11636, nc11637, nc11638, nc11639, nc11640, nc11641, 
        nc11642, nc11643, nc11644, nc11645, \R_DATA_TEMPR7[23] , 
        \R_DATA_TEMPR7[22] }), .B_DOUT({nc11646, nc11647, nc11648, 
        nc11649, nc11650, nc11651, nc11652, nc11653, nc11654, nc11655, 
        nc11656, nc11657, nc11658, nc11659, nc11660, nc11661, nc11662, 
        nc11663, nc11664, nc11665}), .DB_DETECT(\DB_DETECT[7][11] ), 
        .SB_CORRECT(\SB_CORRECT[7][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1 (.A_DOUT({nc11666, 
        nc11667, nc11668, nc11669, nc11670, nc11671, nc11672, nc11673, 
        nc11674, nc11675, nc11676, nc11677, nc11678, nc11679, nc11680, 
        nc11681, nc11682, nc11683, \R_DATA_TEMPR0[3] , 
        \R_DATA_TEMPR0[2] }), .B_DOUT({nc11684, nc11685, nc11686, 
        nc11687, nc11688, nc11689, nc11690, nc11691, nc11692, nc11693, 
        nc11694, nc11695, nc11696, nc11697, nc11698, nc11699, nc11700, 
        nc11701, nc11702, nc11703}), .DB_DETECT(\DB_DETECT[0][1] ), 
        .SB_CORRECT(\SB_CORRECT[0][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C13 (.A_DOUT({
        nc11704, nc11705, nc11706, nc11707, nc11708, nc11709, nc11710, 
        nc11711, nc11712, nc11713, nc11714, nc11715, nc11716, nc11717, 
        nc11718, nc11719, nc11720, nc11721, \R_DATA_TEMPR3[27] , 
        \R_DATA_TEMPR3[26] }), .B_DOUT({nc11722, nc11723, nc11724, 
        nc11725, nc11726, nc11727, nc11728, nc11729, nc11730, nc11731, 
        nc11732, nc11733, nc11734, nc11735, nc11736, nc11737, nc11738, 
        nc11739, nc11740, nc11741}), .DB_DETECT(\DB_DETECT[3][13] ), 
        .SB_CORRECT(\SB_CORRECT[3][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C5 (.A_DOUT({
        nc11742, nc11743, nc11744, nc11745, nc11746, nc11747, nc11748, 
        nc11749, nc11750, nc11751, nc11752, nc11753, nc11754, nc11755, 
        nc11756, nc11757, nc11758, nc11759, \R_DATA_TEMPR26[11] , 
        \R_DATA_TEMPR26[10] }), .B_DOUT({nc11760, nc11761, nc11762, 
        nc11763, nc11764, nc11765, nc11766, nc11767, nc11768, nc11769, 
        nc11770, nc11771, nc11772, nc11773, nc11774, nc11775, nc11776, 
        nc11777, nc11778, nc11779}), .DB_DETECT(\DB_DETECT[26][5] ), 
        .SB_CORRECT(\SB_CORRECT[26][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_84 (.A(OR4_223_Y), .B(OR4_355_Y), .C(OR4_138_Y), .D(
        OR4_291_Y), .Y(OR4_84_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C17 (.A_DOUT({
        nc11780, nc11781, nc11782, nc11783, nc11784, nc11785, nc11786, 
        nc11787, nc11788, nc11789, nc11790, nc11791, nc11792, nc11793, 
        nc11794, nc11795, nc11796, nc11797, \R_DATA_TEMPR27[35] , 
        \R_DATA_TEMPR27[34] }), .B_DOUT({nc11798, nc11799, nc11800, 
        nc11801, nc11802, nc11803, nc11804, nc11805, nc11806, nc11807, 
        nc11808, nc11809, nc11810, nc11811, nc11812, nc11813, nc11814, 
        nc11815, nc11816, nc11817}), .DB_DETECT(\DB_DETECT[27][17] ), 
        .SB_CORRECT(\SB_CORRECT[27][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_148 (.A(\R_DATA_TEMPR12[30] ), .B(\R_DATA_TEMPR13[30] ), 
        .C(\R_DATA_TEMPR14[30] ), .D(\R_DATA_TEMPR15[30] ), .Y(
        OR4_148_Y));
    OR4 OR4_228 (.A(\R_DATA_TEMPR0[18] ), .B(\R_DATA_TEMPR1[18] ), .C(
        \R_DATA_TEMPR2[18] ), .D(\R_DATA_TEMPR3[18] ), .Y(OR4_228_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C18 (.A_DOUT({
        nc11818, nc11819, nc11820, nc11821, nc11822, nc11823, nc11824, 
        nc11825, nc11826, nc11827, nc11828, nc11829, nc11830, nc11831, 
        nc11832, nc11833, nc11834, nc11835, \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR1[36] }), .B_DOUT({nc11836, nc11837, nc11838, 
        nc11839, nc11840, nc11841, nc11842, nc11843, nc11844, nc11845, 
        nc11846, nc11847, nc11848, nc11849, nc11850, nc11851, nc11852, 
        nc11853, nc11854, nc11855}), .DB_DETECT(\DB_DETECT[1][18] ), 
        .SB_CORRECT(\SB_CORRECT[1][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C7 (.A_DOUT({
        nc11856, nc11857, nc11858, nc11859, nc11860, nc11861, nc11862, 
        nc11863, nc11864, nc11865, nc11866, nc11867, nc11868, nc11869, 
        nc11870, nc11871, nc11872, nc11873, \R_DATA_TEMPR30[15] , 
        \R_DATA_TEMPR30[14] }), .B_DOUT({nc11874, nc11875, nc11876, 
        nc11877, nc11878, nc11879, nc11880, nc11881, nc11882, nc11883, 
        nc11884, nc11885, nc11886, nc11887, nc11888, nc11889, nc11890, 
        nc11891, nc11892, nc11893}), .DB_DETECT(\DB_DETECT[30][7] ), 
        .SB_CORRECT(\SB_CORRECT[30][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C19 (.A_DOUT({
        nc11894, nc11895, nc11896, nc11897, nc11898, nc11899, nc11900, 
        nc11901, nc11902, nc11903, nc11904, nc11905, nc11906, nc11907, 
        nc11908, nc11909, nc11910, nc11911, \R_DATA_TEMPR29[39] , 
        \R_DATA_TEMPR29[38] }), .B_DOUT({nc11912, nc11913, nc11914, 
        nc11915, nc11916, nc11917, nc11918, nc11919, nc11920, nc11921, 
        nc11922, nc11923, nc11924, nc11925, nc11926, nc11927, nc11928, 
        nc11929, nc11930, nc11931}), .DB_DETECT(\DB_DETECT[29][19] ), 
        .SB_CORRECT(\SB_CORRECT[29][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C10 (.A_DOUT({
        nc11932, nc11933, nc11934, nc11935, nc11936, nc11937, nc11938, 
        nc11939, nc11940, nc11941, nc11942, nc11943, nc11944, nc11945, 
        nc11946, nc11947, nc11948, nc11949, \R_DATA_TEMPR9[21] , 
        \R_DATA_TEMPR9[20] }), .B_DOUT({nc11950, nc11951, nc11952, 
        nc11953, nc11954, nc11955, nc11956, nc11957, nc11958, nc11959, 
        nc11960, nc11961, nc11962, nc11963, nc11964, nc11965, nc11966, 
        nc11967, nc11968, nc11969}), .DB_DETECT(\DB_DETECT[9][10] ), 
        .SB_CORRECT(\SB_CORRECT[9][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C17 (.A_DOUT({
        nc11970, nc11971, nc11972, nc11973, nc11974, nc11975, nc11976, 
        nc11977, nc11978, nc11979, nc11980, nc11981, nc11982, nc11983, 
        nc11984, nc11985, nc11986, nc11987, \R_DATA_TEMPR0[35] , 
        \R_DATA_TEMPR0[34] }), .B_DOUT({nc11988, nc11989, nc11990, 
        nc11991, nc11992, nc11993, nc11994, nc11995, nc11996, nc11997, 
        nc11998, nc11999, nc12000, nc12001, nc12002, nc12003, nc12004, 
        nc12005, nc12006, nc12007}), .DB_DETECT(\DB_DETECT[0][17] ), 
        .SB_CORRECT(\SB_CORRECT[0][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C8 (.A_DOUT({nc12008, 
        nc12009, nc12010, nc12011, nc12012, nc12013, nc12014, nc12015, 
        nc12016, nc12017, nc12018, nc12019, nc12020, nc12021, nc12022, 
        nc12023, nc12024, nc12025, \R_DATA_TEMPR5[17] , 
        \R_DATA_TEMPR5[16] }), .B_DOUT({nc12026, nc12027, nc12028, 
        nc12029, nc12030, nc12031, nc12032, nc12033, nc12034, nc12035, 
        nc12036, nc12037, nc12038, nc12039, nc12040, nc12041, nc12042, 
        nc12043, nc12044, nc12045}), .DB_DETECT(\DB_DETECT[5][8] ), 
        .SB_CORRECT(\SB_CORRECT[5][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_153 (.A(OR4_184_Y), .B(OR4_19_Y), .C(OR4_159_Y), .D(
        OR4_335_Y), .Y(OR4_153_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C13 (.A_DOUT({
        nc12046, nc12047, nc12048, nc12049, nc12050, nc12051, nc12052, 
        nc12053, nc12054, nc12055, nc12056, nc12057, nc12058, nc12059, 
        nc12060, nc12061, nc12062, nc12063, \R_DATA_TEMPR26[27] , 
        \R_DATA_TEMPR26[26] }), .B_DOUT({nc12064, nc12065, nc12066, 
        nc12067, nc12068, nc12069, nc12070, nc12071, nc12072, nc12073, 
        nc12074, nc12075, nc12076, nc12077, nc12078, nc12079, nc12080, 
        nc12081, nc12082, nc12083}), .DB_DETECT(\DB_DETECT[26][13] ), 
        .SB_CORRECT(\SB_CORRECT[26][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_9 (.A(\R_DATA_TEMPR24[19] ), .B(\R_DATA_TEMPR25[19] ), .C(
        \R_DATA_TEMPR26[19] ), .D(\R_DATA_TEMPR27[19] ), .Y(OR4_9_Y));
    OR4 OR4_231 (.A(\R_DATA_TEMPR0[2] ), .B(\R_DATA_TEMPR1[2] ), .C(
        \R_DATA_TEMPR2[2] ), .D(\R_DATA_TEMPR3[2] ), .Y(OR4_231_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C12 (.A_DOUT({
        nc12084, nc12085, nc12086, nc12087, nc12088, nc12089, nc12090, 
        nc12091, nc12092, nc12093, nc12094, nc12095, nc12096, nc12097, 
        nc12098, nc12099, nc12100, nc12101, \R_DATA_TEMPR31[25] , 
        \R_DATA_TEMPR31[24] }), .B_DOUT({nc12102, nc12103, nc12104, 
        nc12105, nc12106, nc12107, nc12108, nc12109, nc12110, nc12111, 
        nc12112, nc12113, nc12114, nc12115, nc12116, nc12117, nc12118, 
        nc12119, nc12120, nc12121}), .DB_DETECT(\DB_DETECT[31][12] ), 
        .SB_CORRECT(\SB_CORRECT[31][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C3 (.A_DOUT({nc12122, 
        nc12123, nc12124, nc12125, nc12126, nc12127, nc12128, nc12129, 
        nc12130, nc12131, nc12132, nc12133, nc12134, nc12135, nc12136, 
        nc12137, nc12138, nc12139, \R_DATA_TEMPR0[7] , 
        \R_DATA_TEMPR0[6] }), .B_DOUT({nc12140, nc12141, nc12142, 
        nc12143, nc12144, nc12145, nc12146, nc12147, nc12148, nc12149, 
        nc12150, nc12151, nc12152, nc12153, nc12154, nc12155, nc12156, 
        nc12157, nc12158, nc12159}), .DB_DETECT(\DB_DETECT[0][3] ), 
        .SB_CORRECT(\SB_CORRECT[0][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C3 (.A_DOUT({nc12160, 
        nc12161, nc12162, nc12163, nc12164, nc12165, nc12166, nc12167, 
        nc12168, nc12169, nc12170, nc12171, nc12172, nc12173, nc12174, 
        nc12175, nc12176, nc12177, \R_DATA_TEMPR8[7] , 
        \R_DATA_TEMPR8[6] }), .B_DOUT({nc12178, nc12179, nc12180, 
        nc12181, nc12182, nc12183, nc12184, nc12185, nc12186, nc12187, 
        nc12188, nc12189, nc12190, nc12191, nc12192, nc12193, nc12194, 
        nc12195, nc12196, nc12197}), .DB_DETECT(\DB_DETECT[8][3] ), 
        .SB_CORRECT(\SB_CORRECT[8][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C7 (.A_DOUT({
        nc12198, nc12199, nc12200, nc12201, nc12202, nc12203, nc12204, 
        nc12205, nc12206, nc12207, nc12208, nc12209, nc12210, nc12211, 
        nc12212, nc12213, nc12214, nc12215, \R_DATA_TEMPR31[15] , 
        \R_DATA_TEMPR31[14] }), .B_DOUT({nc12216, nc12217, nc12218, 
        nc12219, nc12220, nc12221, nc12222, nc12223, nc12224, nc12225, 
        nc12226, nc12227, nc12228, nc12229, nc12230, nc12231, nc12232, 
        nc12233, nc12234, nc12235}), .DB_DETECT(\DB_DETECT[31][7] ), 
        .SB_CORRECT(\SB_CORRECT[31][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_104 (.A(\R_DATA_TEMPR12[2] ), .B(\R_DATA_TEMPR13[2] ), .C(
        \R_DATA_TEMPR14[2] ), .D(\R_DATA_TEMPR15[2] ), .Y(OR4_104_Y));
    OR4 OR4_292 (.A(OR4_326_Y), .B(OR4_4_Y), .C(OR4_24_Y), .D(OR4_6_Y), 
        .Y(OR4_292_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C11 (.A_DOUT({
        nc12236, nc12237, nc12238, nc12239, nc12240, nc12241, nc12242, 
        nc12243, nc12244, nc12245, nc12246, nc12247, nc12248, nc12249, 
        nc12250, nc12251, nc12252, nc12253, \R_DATA_TEMPR5[23] , 
        \R_DATA_TEMPR5[22] }), .B_DOUT({nc12254, nc12255, nc12256, 
        nc12257, nc12258, nc12259, nc12260, nc12261, nc12262, nc12263, 
        nc12264, nc12265, nc12266, nc12267, nc12268, nc12269, nc12270, 
        nc12271, nc12272, nc12273}), .DB_DETECT(\DB_DETECT[5][11] ), 
        .SB_CORRECT(\SB_CORRECT[5][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C17 (.A_DOUT({
        nc12274, nc12275, nc12276, nc12277, nc12278, nc12279, nc12280, 
        nc12281, nc12282, nc12283, nc12284, nc12285, nc12286, nc12287, 
        nc12288, nc12289, nc12290, nc12291, \R_DATA_TEMPR18[35] , 
        \R_DATA_TEMPR18[34] }), .B_DOUT({nc12292, nc12293, nc12294, 
        nc12295, nc12296, nc12297, nc12298, nc12299, nc12300, nc12301, 
        nc12302, nc12303, nc12304, nc12305, nc12306, nc12307, nc12308, 
        nc12309, nc12310, nc12311}), .DB_DETECT(\DB_DETECT[18][17] ), 
        .SB_CORRECT(\SB_CORRECT[18][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C13 (.A_DOUT({
        nc12312, nc12313, nc12314, nc12315, nc12316, nc12317, nc12318, 
        nc12319, nc12320, nc12321, nc12322, nc12323, nc12324, nc12325, 
        nc12326, nc12327, nc12328, nc12329, \R_DATA_TEMPR12[27] , 
        \R_DATA_TEMPR12[26] }), .B_DOUT({nc12330, nc12331, nc12332, 
        nc12333, nc12334, nc12335, nc12336, nc12337, nc12338, nc12339, 
        nc12340, nc12341, nc12342, nc12343, nc12344, nc12345, nc12346, 
        nc12347, nc12348, nc12349}), .DB_DETECT(\DB_DETECT[12][13] ), 
        .SB_CORRECT(\SB_CORRECT[12][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C19 (.A_DOUT({
        nc12350, nc12351, nc12352, nc12353, nc12354, nc12355, nc12356, 
        nc12357, nc12358, nc12359, nc12360, nc12361, nc12362, nc12363, 
        nc12364, nc12365, nc12366, nc12367, \R_DATA_TEMPR6[39] , 
        \R_DATA_TEMPR6[38] }), .B_DOUT({nc12368, nc12369, nc12370, 
        nc12371, nc12372, nc12373, nc12374, nc12375, nc12376, nc12377, 
        nc12378, nc12379, nc12380, nc12381, nc12382, nc12383, nc12384, 
        nc12385, nc12386, nc12387}), .DB_DETECT(\DB_DETECT[6][19] ), 
        .SB_CORRECT(\SB_CORRECT[6][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_174 (.A(OR4_47_Y), .B(OR4_75_Y), .C(OR4_190_Y), .D(
        OR4_71_Y), .Y(OR4_174_Y));
    OR2 OR2_34 (.A(\R_DATA_TEMPR20[1] ), .B(\R_DATA_TEMPR21[1] ), .Y(
        OR2_34_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C14 (.A_DOUT({
        nc12388, nc12389, nc12390, nc12391, nc12392, nc12393, nc12394, 
        nc12395, nc12396, nc12397, nc12398, nc12399, nc12400, nc12401, 
        nc12402, nc12403, nc12404, nc12405, \R_DATA_TEMPR27[29] , 
        \R_DATA_TEMPR27[28] }), .B_DOUT({nc12406, nc12407, nc12408, 
        nc12409, nc12410, nc12411, nc12412, nc12413, nc12414, nc12415, 
        nc12416, nc12417, nc12418, nc12419, nc12420, nc12421, nc12422, 
        nc12423, nc12424, nc12425}), .DB_DETECT(\DB_DETECT[27][14] ), 
        .SB_CORRECT(\SB_CORRECT[27][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C3 (.A_DOUT({
        nc12426, nc12427, nc12428, nc12429, nc12430, nc12431, nc12432, 
        nc12433, nc12434, nc12435, nc12436, nc12437, nc12438, nc12439, 
        nc12440, nc12441, nc12442, nc12443, \R_DATA_TEMPR22[7] , 
        \R_DATA_TEMPR22[6] }), .B_DOUT({nc12444, nc12445, nc12446, 
        nc12447, nc12448, nc12449, nc12450, nc12451, nc12452, nc12453, 
        nc12454, nc12455, nc12456, nc12457, nc12458, nc12459, nc12460, 
        nc12461, nc12462, nc12463}), .DB_DETECT(\DB_DETECT[22][3] ), 
        .SB_CORRECT(\SB_CORRECT[22][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C6 (.A_DOUT({
        nc12464, nc12465, nc12466, nc12467, nc12468, nc12469, nc12470, 
        nc12471, nc12472, nc12473, nc12474, nc12475, nc12476, nc12477, 
        nc12478, nc12479, nc12480, nc12481, \R_DATA_TEMPR13[13] , 
        \R_DATA_TEMPR13[12] }), .B_DOUT({nc12482, nc12483, nc12484, 
        nc12485, nc12486, nc12487, nc12488, nc12489, nc12490, nc12491, 
        nc12492, nc12493, nc12494, nc12495, nc12496, nc12497, nc12498, 
        nc12499, nc12500, nc12501}), .DB_DETECT(\DB_DETECT[13][6] ), 
        .SB_CORRECT(\SB_CORRECT[13][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_56 (.A(\R_DATA_TEMPR24[37] ), .B(\R_DATA_TEMPR25[37] ), .C(
        \R_DATA_TEMPR26[37] ), .D(\R_DATA_TEMPR27[37] ), .Y(OR4_56_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0 (.A_DOUT({nc12502, 
        nc12503, nc12504, nc12505, nc12506, nc12507, nc12508, nc12509, 
        nc12510, nc12511, nc12512, nc12513, nc12514, nc12515, nc12516, 
        nc12517, nc12518, nc12519, \R_DATA_TEMPR5[1] , 
        \R_DATA_TEMPR5[0] }), .B_DOUT({nc12520, nc12521, nc12522, 
        nc12523, nc12524, nc12525, nc12526, nc12527, nc12528, nc12529, 
        nc12530, nc12531, nc12532, nc12533, nc12534, nc12535, nc12536, 
        nc12537, nc12538, nc12539}), .DB_DETECT(\DB_DETECT[5][0] ), 
        .SB_CORRECT(\SB_CORRECT[5][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0 (.A_DOUT({
        nc12540, nc12541, nc12542, nc12543, nc12544, nc12545, nc12546, 
        nc12547, nc12548, nc12549, nc12550, nc12551, nc12552, nc12553, 
        nc12554, nc12555, nc12556, nc12557, \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR12[0] }), .B_DOUT({nc12558, nc12559, nc12560, 
        nc12561, nc12562, nc12563, nc12564, nc12565, nc12566, nc12567, 
        nc12568, nc12569, nc12570, nc12571, nc12572, nc12573, nc12574, 
        nc12575, nc12576, nc12577}), .DB_DETECT(\DB_DETECT[12][0] ), 
        .SB_CORRECT(\SB_CORRECT[12][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C7 (.A_DOUT({nc12578, 
        nc12579, nc12580, nc12581, nc12582, nc12583, nc12584, nc12585, 
        nc12586, nc12587, nc12588, nc12589, nc12590, nc12591, nc12592, 
        nc12593, nc12594, nc12595, \R_DATA_TEMPR6[15] , 
        \R_DATA_TEMPR6[14] }), .B_DOUT({nc12596, nc12597, nc12598, 
        nc12599, nc12600, nc12601, nc12602, nc12603, nc12604, nc12605, 
        nc12606, nc12607, nc12608, nc12609, nc12610, nc12611, nc12612, 
        nc12613, nc12614, nc12615}), .DB_DETECT(\DB_DETECT[6][7] ), 
        .SB_CORRECT(\SB_CORRECT[6][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[2]  (.A(CFG2_1_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[2] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C18 (.A_DOUT({
        nc12616, nc12617, nc12618, nc12619, nc12620, nc12621, nc12622, 
        nc12623, nc12624, nc12625, nc12626, nc12627, nc12628, nc12629, 
        nc12630, nc12631, nc12632, nc12633, \R_DATA_TEMPR29[37] , 
        \R_DATA_TEMPR29[36] }), .B_DOUT({nc12634, nc12635, nc12636, 
        nc12637, nc12638, nc12639, nc12640, nc12641, nc12642, nc12643, 
        nc12644, nc12645, nc12646, nc12647, nc12648, nc12649, nc12650, 
        nc12651, nc12652, nc12653}), .DB_DETECT(\DB_DETECT[29][18] ), 
        .SB_CORRECT(\SB_CORRECT[29][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[2]  (.A(OR4_192_Y), .B(OR4_170_Y), .C(OR4_243_Y), 
        .D(OR4_274_Y), .Y(R_DATA[2]));
    OR4 OR4_152 (.A(\R_DATA_TEMPR28[24] ), .B(\R_DATA_TEMPR29[24] ), 
        .C(\R_DATA_TEMPR30[24] ), .D(\R_DATA_TEMPR31[24] ), .Y(
        OR4_152_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C5 (.A_DOUT({
        nc12654, nc12655, nc12656, nc12657, nc12658, nc12659, nc12660, 
        nc12661, nc12662, nc12663, nc12664, nc12665, nc12666, nc12667, 
        nc12668, nc12669, nc12670, nc12671, \R_DATA_TEMPR18[11] , 
        \R_DATA_TEMPR18[10] }), .B_DOUT({nc12672, nc12673, nc12674, 
        nc12675, nc12676, nc12677, nc12678, nc12679, nc12680, nc12681, 
        nc12682, nc12683, nc12684, nc12685, nc12686, nc12687, nc12688, 
        nc12689, nc12690, nc12691}), .DB_DETECT(\DB_DETECT[18][5] ), 
        .SB_CORRECT(\SB_CORRECT[18][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C17 (.A_DOUT({
        nc12692, nc12693, nc12694, nc12695, nc12696, nc12697, nc12698, 
        nc12699, nc12700, nc12701, nc12702, nc12703, nc12704, nc12705, 
        nc12706, nc12707, nc12708, nc12709, \R_DATA_TEMPR22[35] , 
        \R_DATA_TEMPR22[34] }), .B_DOUT({nc12710, nc12711, nc12712, 
        nc12713, nc12714, nc12715, nc12716, nc12717, nc12718, nc12719, 
        nc12720, nc12721, nc12722, nc12723, nc12724, nc12725, nc12726, 
        nc12727, nc12728, nc12729}), .DB_DETECT(\DB_DETECT[22][17] ), 
        .SB_CORRECT(\SB_CORRECT[22][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C18 (.A_DOUT({
        nc12730, nc12731, nc12732, nc12733, nc12734, nc12735, nc12736, 
        nc12737, nc12738, nc12739, nc12740, nc12741, nc12742, nc12743, 
        nc12744, nc12745, nc12746, nc12747, \R_DATA_TEMPR8[37] , 
        \R_DATA_TEMPR8[36] }), .B_DOUT({nc12748, nc12749, nc12750, 
        nc12751, nc12752, nc12753, nc12754, nc12755, nc12756, nc12757, 
        nc12758, nc12759, nc12760, nc12761, nc12762, nc12763, nc12764, 
        nc12765, nc12766, nc12767}), .DB_DETECT(\DB_DETECT[8][18] ), 
        .SB_CORRECT(\SB_CORRECT[8][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_39 (.A(\R_DATA_TEMPR8[4] ), .B(\R_DATA_TEMPR9[4] ), .C(
        \R_DATA_TEMPR10[4] ), .D(\R_DATA_TEMPR11[4] ), .Y(OR4_39_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C16 (.A_DOUT({
        nc12768, nc12769, nc12770, nc12771, nc12772, nc12773, nc12774, 
        nc12775, nc12776, nc12777, nc12778, nc12779, nc12780, nc12781, 
        nc12782, nc12783, nc12784, nc12785, \R_DATA_TEMPR26[33] , 
        \R_DATA_TEMPR26[32] }), .B_DOUT({nc12786, nc12787, nc12788, 
        nc12789, nc12790, nc12791, nc12792, nc12793, nc12794, nc12795, 
        nc12796, nc12797, nc12798, nc12799, nc12800, nc12801, nc12802, 
        nc12803, nc12804, nc12805}), .DB_DETECT(\DB_DETECT[26][16] ), 
        .SB_CORRECT(\SB_CORRECT[26][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_211 (.A(OR4_161_Y), .B(OR2_36_Y), .C(\R_DATA_TEMPR22[27] ), 
        .D(\R_DATA_TEMPR23[27] ), .Y(OR4_211_Y));
    OR2 OR2_9 (.A(\R_DATA_TEMPR20[3] ), .B(\R_DATA_TEMPR21[3] ), .Y(
        OR2_9_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C19 (.A_DOUT({
        nc12806, nc12807, nc12808, nc12809, nc12810, nc12811, nc12812, 
        nc12813, nc12814, nc12815, nc12816, nc12817, nc12818, nc12819, 
        nc12820, nc12821, nc12822, nc12823, \R_DATA_TEMPR13[39] , 
        \R_DATA_TEMPR13[38] }), .B_DOUT({nc12824, nc12825, nc12826, 
        nc12827, nc12828, nc12829, nc12830, nc12831, nc12832, nc12833, 
        nc12834, nc12835, nc12836, nc12837, nc12838, nc12839, nc12840, 
        nc12841, nc12842, nc12843}), .DB_DETECT(\DB_DETECT[13][19] ), 
        .SB_CORRECT(\SB_CORRECT[13][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C8 (.A_DOUT({nc12844, 
        nc12845, nc12846, nc12847, nc12848, nc12849, nc12850, nc12851, 
        nc12852, nc12853, nc12854, nc12855, nc12856, nc12857, nc12858, 
        nc12859, nc12860, nc12861, \R_DATA_TEMPR6[17] , 
        \R_DATA_TEMPR6[16] }), .B_DOUT({nc12862, nc12863, nc12864, 
        nc12865, nc12866, nc12867, nc12868, nc12869, nc12870, nc12871, 
        nc12872, nc12873, nc12874, nc12875, nc12876, nc12877, nc12878, 
        nc12879, nc12880, nc12881}), .DB_DETECT(\DB_DETECT[6][8] ), 
        .SB_CORRECT(\SB_CORRECT[6][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C5 (.A_DOUT({
        nc12882, nc12883, nc12884, nc12885, nc12886, nc12887, nc12888, 
        nc12889, nc12890, nc12891, nc12892, nc12893, nc12894, nc12895, 
        nc12896, nc12897, nc12898, nc12899, \R_DATA_TEMPR21[11] , 
        \R_DATA_TEMPR21[10] }), .B_DOUT({nc12900, nc12901, nc12902, 
        nc12903, nc12904, nc12905, nc12906, nc12907, nc12908, nc12909, 
        nc12910, nc12911, nc12912, nc12913, nc12914, nc12915, nc12916, 
        nc12917, nc12918, nc12919}), .DB_DETECT(\DB_DETECT[21][5] ), 
        .SB_CORRECT(\SB_CORRECT[21][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[21][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_222 (.A(\R_DATA_TEMPR24[5] ), .B(\R_DATA_TEMPR25[5] ), .C(
        \R_DATA_TEMPR26[5] ), .D(\R_DATA_TEMPR27[5] ), .Y(OR4_222_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C5 (.A_DOUT({
        nc12920, nc12921, nc12922, nc12923, nc12924, nc12925, nc12926, 
        nc12927, nc12928, nc12929, nc12930, nc12931, nc12932, nc12933, 
        nc12934, nc12935, nc12936, nc12937, \R_DATA_TEMPR24[11] , 
        \R_DATA_TEMPR24[10] }), .B_DOUT({nc12938, nc12939, nc12940, 
        nc12941, nc12942, nc12943, nc12944, nc12945, nc12946, nc12947, 
        nc12948, nc12949, nc12950, nc12951, nc12952, nc12953, nc12954, 
        nc12955, nc12956, nc12957}), .DB_DETECT(\DB_DETECT[24][5] ), 
        .SB_CORRECT(\SB_CORRECT[24][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_145 (.A(\R_DATA_TEMPR8[21] ), .B(\R_DATA_TEMPR9[21] ), .C(
        \R_DATA_TEMPR10[21] ), .D(\R_DATA_TEMPR11[21] ), .Y(OR4_145_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C15 (.A_DOUT({
        nc12958, nc12959, nc12960, nc12961, nc12962, nc12963, nc12964, 
        nc12965, nc12966, nc12967, nc12968, nc12969, nc12970, nc12971, 
        nc12972, nc12973, nc12974, nc12975, \R_DATA_TEMPR26[31] , 
        \R_DATA_TEMPR26[30] }), .B_DOUT({nc12976, nc12977, nc12978, 
        nc12979, nc12980, nc12981, nc12982, nc12983, nc12984, nc12985, 
        nc12986, nc12987, nc12988, nc12989, nc12990, nc12991, nc12992, 
        nc12993, nc12994, nc12995}), .DB_DETECT(\DB_DETECT[26][15] ), 
        .SB_CORRECT(\SB_CORRECT[26][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C3 (.A_DOUT({nc12996, 
        nc12997, nc12998, nc12999, nc13000, nc13001, nc13002, nc13003, 
        nc13004, nc13005, nc13006, nc13007, nc13008, nc13009, nc13010, 
        nc13011, nc13012, nc13013, \R_DATA_TEMPR2[7] , 
        \R_DATA_TEMPR2[6] }), .B_DOUT({nc13014, nc13015, nc13016, 
        nc13017, nc13018, nc13019, nc13020, nc13021, nc13022, nc13023, 
        nc13024, nc13025, nc13026, nc13027, nc13028, nc13029, nc13030, 
        nc13031, nc13032, nc13033}), .DB_DETECT(\DB_DETECT[2][3] ), 
        .SB_CORRECT(\SB_CORRECT[2][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C4 (.A_DOUT({nc13034, 
        nc13035, nc13036, nc13037, nc13038, nc13039, nc13040, nc13041, 
        nc13042, nc13043, nc13044, nc13045, nc13046, nc13047, nc13048, 
        nc13049, nc13050, nc13051, \R_DATA_TEMPR4[9] , 
        \R_DATA_TEMPR4[8] }), .B_DOUT({nc13052, nc13053, nc13054, 
        nc13055, nc13056, nc13057, nc13058, nc13059, nc13060, nc13061, 
        nc13062, nc13063, nc13064, nc13065, nc13066, nc13067, nc13068, 
        nc13069, nc13070, nc13071}), .DB_DETECT(\DB_DETECT[4][4] ), 
        .SB_CORRECT(\SB_CORRECT[4][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_16 (.A(\R_DATA_TEMPR4[19] ), .B(\R_DATA_TEMPR5[19] ), .C(
        \R_DATA_TEMPR6[19] ), .D(\R_DATA_TEMPR7[19] ), .Y(OR4_16_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C4 (.A_DOUT({nc13072, 
        nc13073, nc13074, nc13075, nc13076, nc13077, nc13078, nc13079, 
        nc13080, nc13081, nc13082, nc13083, nc13084, nc13085, nc13086, 
        nc13087, nc13088, nc13089, \R_DATA_TEMPR3[9] , 
        \R_DATA_TEMPR3[8] }), .B_DOUT({nc13090, nc13091, nc13092, 
        nc13093, nc13094, nc13095, nc13096, nc13097, nc13098, nc13099, 
        nc13100, nc13101, nc13102, nc13103, nc13104, nc13105, nc13106, 
        nc13107, nc13108, nc13109}), .DB_DETECT(\DB_DETECT[3][4] ), 
        .SB_CORRECT(\SB_CORRECT[3][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_259 (.A(\R_DATA_TEMPR24[30] ), .B(\R_DATA_TEMPR25[30] ), 
        .C(\R_DATA_TEMPR26[30] ), .D(\R_DATA_TEMPR27[30] ), .Y(
        OR4_259_Y));
    OR4 OR4_331 (.A(OR4_49_Y), .B(OR2_2_Y), .C(\R_DATA_TEMPR22[26] ), 
        .D(\R_DATA_TEMPR23[26] ), .Y(OR4_331_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C8 (.A_DOUT({
        nc13110, nc13111, nc13112, nc13113, nc13114, nc13115, nc13116, 
        nc13117, nc13118, nc13119, nc13120, nc13121, nc13122, nc13123, 
        nc13124, nc13125, nc13126, nc13127, \R_DATA_TEMPR22[17] , 
        \R_DATA_TEMPR22[16] }), .B_DOUT({nc13128, nc13129, nc13130, 
        nc13131, nc13132, nc13133, nc13134, nc13135, nc13136, nc13137, 
        nc13138, nc13139, nc13140, nc13141, nc13142, nc13143, nc13144, 
        nc13145, nc13146, nc13147}), .DB_DETECT(\DB_DETECT[22][8] ), 
        .SB_CORRECT(\SB_CORRECT[22][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_4 (.A(\R_DATA_TEMPR4[1] ), .B(\R_DATA_TEMPR5[1] ), .C(
        \R_DATA_TEMPR6[1] ), .D(\R_DATA_TEMPR7[1] ), .Y(OR4_4_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C6 (.A_DOUT({nc13148, 
        nc13149, nc13150, nc13151, nc13152, nc13153, nc13154, nc13155, 
        nc13156, nc13157, nc13158, nc13159, nc13160, nc13161, nc13162, 
        nc13163, nc13164, nc13165, \R_DATA_TEMPR1[13] , 
        \R_DATA_TEMPR1[12] }), .B_DOUT({nc13166, nc13167, nc13168, 
        nc13169, nc13170, nc13171, nc13172, nc13173, nc13174, nc13175, 
        nc13176, nc13177, nc13178, nc13179, nc13180, nc13181, nc13182, 
        nc13183, nc13184, nc13185}), .DB_DETECT(\DB_DETECT[1][6] ), 
        .SB_CORRECT(\SB_CORRECT[1][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_320 (.A(\R_DATA_TEMPR24[21] ), .B(\R_DATA_TEMPR25[21] ), 
        .C(\R_DATA_TEMPR26[21] ), .D(\R_DATA_TEMPR27[21] ), .Y(
        OR4_320_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C14 (.A_DOUT({
        nc13186, nc13187, nc13188, nc13189, nc13190, nc13191, nc13192, 
        nc13193, nc13194, nc13195, nc13196, nc13197, nc13198, nc13199, 
        nc13200, nc13201, nc13202, nc13203, \R_DATA_TEMPR22[29] , 
        \R_DATA_TEMPR22[28] }), .B_DOUT({nc13204, nc13205, nc13206, 
        nc13207, nc13208, nc13209, nc13210, nc13211, nc13212, nc13213, 
        nc13214, nc13215, nc13216, nc13217, nc13218, nc13219, nc13220, 
        nc13221, nc13222, nc13223}), .DB_DETECT(\DB_DETECT[22][14] ), 
        .SB_CORRECT(\SB_CORRECT[22][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C8 (.A_DOUT({nc13224, 
        nc13225, nc13226, nc13227, nc13228, nc13229, nc13230, nc13231, 
        nc13232, nc13233, nc13234, nc13235, nc13236, nc13237, nc13238, 
        nc13239, nc13240, nc13241, \R_DATA_TEMPR9[17] , 
        \R_DATA_TEMPR9[16] }), .B_DOUT({nc13242, nc13243, nc13244, 
        nc13245, nc13246, nc13247, nc13248, nc13249, nc13250, nc13251, 
        nc13252, nc13253, nc13254, nc13255, nc13256, nc13257, nc13258, 
        nc13259, nc13260, nc13261}), .DB_DETECT(\DB_DETECT[9][8] ), 
        .SB_CORRECT(\SB_CORRECT[9][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[14]  (.A(OR4_342_Y), .B(OR4_210_Y), .C(OR4_23_Y), 
        .D(OR4_185_Y), .Y(R_DATA[14]));
    OR4 OR4_245 (.A(OR4_100_Y), .B(OR2_0_Y), .C(\R_DATA_TEMPR22[12] ), 
        .D(\R_DATA_TEMPR23[12] ), .Y(OR4_245_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C12 (.A_DOUT({
        nc13262, nc13263, nc13264, nc13265, nc13266, nc13267, nc13268, 
        nc13269, nc13270, nc13271, nc13272, nc13273, nc13274, nc13275, 
        nc13276, nc13277, nc13278, nc13279, \R_DATA_TEMPR29[25] , 
        \R_DATA_TEMPR29[24] }), .B_DOUT({nc13280, nc13281, nc13282, 
        nc13283, nc13284, nc13285, nc13286, nc13287, nc13288, nc13289, 
        nc13290, nc13291, nc13292, nc13293, nc13294, nc13295, nc13296, 
        nc13297, nc13298, nc13299}), .DB_DETECT(\DB_DETECT[29][12] ), 
        .SB_CORRECT(\SB_CORRECT[29][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C15 (.A_DOUT({
        nc13300, nc13301, nc13302, nc13303, nc13304, nc13305, nc13306, 
        nc13307, nc13308, nc13309, nc13310, nc13311, nc13312, nc13313, 
        nc13314, nc13315, nc13316, nc13317, \R_DATA_TEMPR2[31] , 
        \R_DATA_TEMPR2[30] }), .B_DOUT({nc13318, nc13319, nc13320, 
        nc13321, nc13322, nc13323, nc13324, nc13325, nc13326, nc13327, 
        nc13328, nc13329, nc13330, nc13331, nc13332, nc13333, nc13334, 
        nc13335, nc13336, nc13337}), .DB_DETECT(\DB_DETECT[2][15] ), 
        .SB_CORRECT(\SB_CORRECT[2][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C10 (.A_DOUT({
        nc13338, nc13339, nc13340, nc13341, nc13342, nc13343, nc13344, 
        nc13345, nc13346, nc13347, nc13348, nc13349, nc13350, nc13351, 
        nc13352, nc13353, nc13354, nc13355, \R_DATA_TEMPR29[21] , 
        \R_DATA_TEMPR29[20] }), .B_DOUT({nc13356, nc13357, nc13358, 
        nc13359, nc13360, nc13361, nc13362, nc13363, nc13364, nc13365, 
        nc13366, nc13367, nc13368, nc13369, nc13370, nc13371, nc13372, 
        nc13373, nc13374, nc13375}), .DB_DETECT(\DB_DETECT[29][10] ), 
        .SB_CORRECT(\SB_CORRECT[29][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_50 (.A(\R_DATA_TEMPR16[5] ), .B(\R_DATA_TEMPR17[5] ), .C(
        \R_DATA_TEMPR18[5] ), .D(\R_DATA_TEMPR19[5] ), .Y(OR4_50_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C13 (.A_DOUT({
        nc13376, nc13377, nc13378, nc13379, nc13380, nc13381, nc13382, 
        nc13383, nc13384, nc13385, nc13386, nc13387, nc13388, nc13389, 
        nc13390, nc13391, nc13392, nc13393, \R_DATA_TEMPR0[27] , 
        \R_DATA_TEMPR0[26] }), .B_DOUT({nc13394, nc13395, nc13396, 
        nc13397, nc13398, nc13399, nc13400, nc13401, nc13402, nc13403, 
        nc13404, nc13405, nc13406, nc13407, nc13408, nc13409, nc13410, 
        nc13411, nc13412, nc13413}), .DB_DETECT(\DB_DETECT[0][13] ), 
        .SB_CORRECT(\SB_CORRECT[0][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_57 (.A(\R_DATA_TEMPR0[36] ), .B(\R_DATA_TEMPR1[36] ), .C(
        \R_DATA_TEMPR2[36] ), .D(\R_DATA_TEMPR3[36] ), .Y(OR4_57_Y));
    OR4 OR4_32 (.A(\R_DATA_TEMPR16[20] ), .B(\R_DATA_TEMPR17[20] ), .C(
        \R_DATA_TEMPR18[20] ), .D(\R_DATA_TEMPR19[20] ), .Y(OR4_32_Y));
    OR4 OR4_260 (.A(\R_DATA_TEMPR28[38] ), .B(\R_DATA_TEMPR29[38] ), 
        .C(\R_DATA_TEMPR30[38] ), .D(\R_DATA_TEMPR31[38] ), .Y(
        OR4_260_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C13 (.A_DOUT({
        nc13414, nc13415, nc13416, nc13417, nc13418, nc13419, nc13420, 
        nc13421, nc13422, nc13423, nc13424, nc13425, nc13426, nc13427, 
        nc13428, nc13429, nc13430, nc13431, \R_DATA_TEMPR27[27] , 
        \R_DATA_TEMPR27[26] }), .B_DOUT({nc13432, nc13433, nc13434, 
        nc13435, nc13436, nc13437, nc13438, nc13439, nc13440, nc13441, 
        nc13442, nc13443, nc13444, nc13445, nc13446, nc13447, nc13448, 
        nc13449, nc13450, nc13451}), .DB_DETECT(\DB_DETECT[27][13] ), 
        .SB_CORRECT(\SB_CORRECT[27][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0 (.A_DOUT({
        nc13452, nc13453, nc13454, nc13455, nc13456, nc13457, nc13458, 
        nc13459, nc13460, nc13461, nc13462, nc13463, nc13464, nc13465, 
        nc13466, nc13467, nc13468, nc13469, \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR30[0] }), .B_DOUT({nc13470, nc13471, nc13472, 
        nc13473, nc13474, nc13475, nc13476, nc13477, nc13478, nc13479, 
        nc13480, nc13481, nc13482, nc13483, nc13484, nc13485, nc13486, 
        nc13487, nc13488, nc13489}), .DB_DETECT(\DB_DETECT[30][0] ), 
        .SB_CORRECT(\SB_CORRECT[30][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C16 (.A_DOUT({
        nc13490, nc13491, nc13492, nc13493, nc13494, nc13495, nc13496, 
        nc13497, nc13498, nc13499, nc13500, nc13501, nc13502, nc13503, 
        nc13504, nc13505, nc13506, nc13507, \R_DATA_TEMPR19[33] , 
        \R_DATA_TEMPR19[32] }), .B_DOUT({nc13508, nc13509, nc13510, 
        nc13511, nc13512, nc13513, nc13514, nc13515, nc13516, nc13517, 
        nc13518, nc13519, nc13520, nc13521, nc13522, nc13523, nc13524, 
        nc13525, nc13526, nc13527}), .DB_DETECT(\DB_DETECT[19][16] ), 
        .SB_CORRECT(\SB_CORRECT[19][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C1 (.A_DOUT({
        nc13528, nc13529, nc13530, nc13531, nc13532, nc13533, nc13534, 
        nc13535, nc13536, nc13537, nc13538, nc13539, nc13540, nc13541, 
        nc13542, nc13543, nc13544, nc13545, \R_DATA_TEMPR23[3] , 
        \R_DATA_TEMPR23[2] }), .B_DOUT({nc13546, nc13547, nc13548, 
        nc13549, nc13550, nc13551, nc13552, nc13553, nc13554, nc13555, 
        nc13556, nc13557, nc13558, nc13559, nc13560, nc13561, nc13562, 
        nc13563, nc13564, nc13565}), .DB_DETECT(\DB_DETECT[23][1] ), 
        .SB_CORRECT(\SB_CORRECT[23][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C15 (.A_DOUT({
        nc13566, nc13567, nc13568, nc13569, nc13570, nc13571, nc13572, 
        nc13573, nc13574, nc13575, nc13576, nc13577, nc13578, nc13579, 
        nc13580, nc13581, nc13582, nc13583, \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR7[30] }), .B_DOUT({nc13584, nc13585, nc13586, 
        nc13587, nc13588, nc13589, nc13590, nc13591, nc13592, nc13593, 
        nc13594, nc13595, nc13596, nc13597, nc13598, nc13599, nc13600, 
        nc13601, nc13602, nc13603}), .DB_DETECT(\DB_DETECT[7][15] ), 
        .SB_CORRECT(\SB_CORRECT[7][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_311 (.A(OR4_52_Y), .B(OR2_29_Y), .C(\R_DATA_TEMPR22[21] ), 
        .D(\R_DATA_TEMPR23[21] ), .Y(OR4_311_Y));
    OR4 OR4_184 (.A(\R_DATA_TEMPR0[37] ), .B(\R_DATA_TEMPR1[37] ), .C(
        \R_DATA_TEMPR2[37] ), .D(\R_DATA_TEMPR3[37] ), .Y(OR4_184_Y));
    OR4 OR4_248 (.A(\R_DATA_TEMPR8[16] ), .B(\R_DATA_TEMPR9[16] ), .C(
        \R_DATA_TEMPR10[16] ), .D(\R_DATA_TEMPR11[16] ), .Y(OR4_248_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C9 (.A_DOUT({nc13604, 
        nc13605, nc13606, nc13607, nc13608, nc13609, nc13610, nc13611, 
        nc13612, nc13613, nc13614, nc13615, nc13616, nc13617, nc13618, 
        nc13619, nc13620, nc13621, \R_DATA_TEMPR7[19] , 
        \R_DATA_TEMPR7[18] }), .B_DOUT({nc13622, nc13623, nc13624, 
        nc13625, nc13626, nc13627, nc13628, nc13629, nc13630, nc13631, 
        nc13632, nc13633, nc13634, nc13635, nc13636, nc13637, nc13638, 
        nc13639, nc13640, nc13641}), .DB_DETECT(\DB_DETECT[7][9] ), 
        .SB_CORRECT(\SB_CORRECT[7][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C5 (.A_DOUT({
        nc13642, nc13643, nc13644, nc13645, nc13646, nc13647, nc13648, 
        nc13649, nc13650, nc13651, nc13652, nc13653, nc13654, nc13655, 
        nc13656, nc13657, nc13658, nc13659, \R_DATA_TEMPR10[11] , 
        \R_DATA_TEMPR10[10] }), .B_DOUT({nc13660, nc13661, nc13662, 
        nc13663, nc13664, nc13665, nc13666, nc13667, nc13668, nc13669, 
        nc13670, nc13671, nc13672, nc13673, nc13674, nc13675, nc13676, 
        nc13677, nc13678, nc13679}), .DB_DETECT(\DB_DETECT[10][5] ), 
        .SB_CORRECT(\SB_CORRECT[10][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0 (.A_DOUT({
        nc13680, nc13681, nc13682, nc13683, nc13684, nc13685, nc13686, 
        nc13687, nc13688, nc13689, nc13690, nc13691, nc13692, nc13693, 
        nc13694, nc13695, nc13696, nc13697, \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR27[0] }), .B_DOUT({nc13698, nc13699, nc13700, 
        nc13701, nc13702, nc13703, nc13704, nc13705, nc13706, nc13707, 
        nc13708, nc13709, nc13710, nc13711, nc13712, nc13713, nc13714, 
        nc13715, nc13716, nc13717}), .DB_DETECT(\DB_DETECT[27][0] ), 
        .SB_CORRECT(\SB_CORRECT[27][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_302 (.A(\R_DATA_TEMPR4[15] ), .B(\R_DATA_TEMPR5[15] ), .C(
        \R_DATA_TEMPR6[15] ), .D(\R_DATA_TEMPR7[15] ), .Y(OR4_302_Y));
    OR4 OR4_266 (.A(\R_DATA_TEMPR0[10] ), .B(\R_DATA_TEMPR1[10] ), .C(
        \R_DATA_TEMPR2[10] ), .D(\R_DATA_TEMPR3[10] ), .Y(OR4_266_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C7 (.A_DOUT({
        nc13718, nc13719, nc13720, nc13721, nc13722, nc13723, nc13724, 
        nc13725, nc13726, nc13727, nc13728, nc13729, nc13730, nc13731, 
        nc13732, nc13733, nc13734, nc13735, \R_DATA_TEMPR23[15] , 
        \R_DATA_TEMPR23[14] }), .B_DOUT({nc13736, nc13737, nc13738, 
        nc13739, nc13740, nc13741, nc13742, nc13743, nc13744, nc13745, 
        nc13746, nc13747, nc13748, nc13749, nc13750, nc13751, nc13752, 
        nc13753, nc13754, nc13755}), .DB_DETECT(\DB_DETECT[23][7] ), 
        .SB_CORRECT(\SB_CORRECT[23][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C16 (.A_DOUT({
        nc13756, nc13757, nc13758, nc13759, nc13760, nc13761, nc13762, 
        nc13763, nc13764, nc13765, nc13766, nc13767, nc13768, nc13769, 
        nc13770, nc13771, nc13772, nc13773, \R_DATA_TEMPR30[33] , 
        \R_DATA_TEMPR30[32] }), .B_DOUT({nc13774, nc13775, nc13776, 
        nc13777, nc13778, nc13779, nc13780, nc13781, nc13782, nc13783, 
        nc13784, nc13785, nc13786, nc13787, nc13788, nc13789, nc13790, 
        nc13791, nc13792, nc13793}), .DB_DETECT(\DB_DETECT[30][16] ), 
        .SB_CORRECT(\SB_CORRECT[30][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_10 (.A(\R_DATA_TEMPR28[20] ), .B(\R_DATA_TEMPR29[20] ), .C(
        \R_DATA_TEMPR30[20] ), .D(\R_DATA_TEMPR31[20] ), .Y(OR4_10_Y));
    OR4 OR4_25 (.A(\R_DATA_TEMPR16[34] ), .B(\R_DATA_TEMPR17[34] ), .C(
        \R_DATA_TEMPR18[34] ), .D(\R_DATA_TEMPR19[34] ), .Y(OR4_25_Y));
    OR4 OR4_76 (.A(\R_DATA_TEMPR0[27] ), .B(\R_DATA_TEMPR1[27] ), .C(
        \R_DATA_TEMPR2[27] ), .D(\R_DATA_TEMPR3[27] ), .Y(OR4_76_Y));
    OR4 OR4_339 (.A(\R_DATA_TEMPR24[17] ), .B(\R_DATA_TEMPR25[17] ), 
        .C(\R_DATA_TEMPR26[17] ), .D(\R_DATA_TEMPR27[17] ), .Y(
        OR4_339_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[4]  (.A(CFG2_4_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[4] ));
    OR4 OR4_193 (.A(OR4_341_Y), .B(OR4_107_Y), .C(OR4_253_Y), .D(
        OR4_38_Y), .Y(OR4_193_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C4 (.A_DOUT({
        nc13794, nc13795, nc13796, nc13797, nc13798, nc13799, nc13800, 
        nc13801, nc13802, nc13803, nc13804, nc13805, nc13806, nc13807, 
        nc13808, nc13809, nc13810, nc13811, \R_DATA_TEMPR30[9] , 
        \R_DATA_TEMPR30[8] }), .B_DOUT({nc13812, nc13813, nc13814, 
        nc13815, nc13816, nc13817, nc13818, nc13819, nc13820, nc13821, 
        nc13822, nc13823, nc13824, nc13825, nc13826, nc13827, nc13828, 
        nc13829, nc13830, nc13831}), .DB_DETECT(\DB_DETECT[30][4] ), 
        .SB_CORRECT(\SB_CORRECT[30][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C12 (.A_DOUT({
        nc13832, nc13833, nc13834, nc13835, nc13836, nc13837, nc13838, 
        nc13839, nc13840, nc13841, nc13842, nc13843, nc13844, nc13845, 
        nc13846, nc13847, nc13848, nc13849, \R_DATA_TEMPR18[25] , 
        \R_DATA_TEMPR18[24] }), .B_DOUT({nc13850, nc13851, nc13852, 
        nc13853, nc13854, nc13855, nc13856, nc13857, nc13858, nc13859, 
        nc13860, nc13861, nc13862, nc13863, nc13864, nc13865, nc13866, 
        nc13867, nc13868, nc13869}), .DB_DETECT(\DB_DETECT[18][12] ), 
        .SB_CORRECT(\SB_CORRECT[18][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C11 (.A_DOUT({
        nc13870, nc13871, nc13872, nc13873, nc13874, nc13875, nc13876, 
        nc13877, nc13878, nc13879, nc13880, nc13881, nc13882, nc13883, 
        nc13884, nc13885, nc13886, nc13887, \R_DATA_TEMPR28[23] , 
        \R_DATA_TEMPR28[22] }), .B_DOUT({nc13888, nc13889, nc13890, 
        nc13891, nc13892, nc13893, nc13894, nc13895, nc13896, nc13897, 
        nc13898, nc13899, nc13900, nc13901, nc13902, nc13903, nc13904, 
        nc13905, nc13906, nc13907}), .DB_DETECT(\DB_DETECT[28][11] ), 
        .SB_CORRECT(\SB_CORRECT[28][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[28][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_17 (.A(\R_DATA_TEMPR12[34] ), .B(\R_DATA_TEMPR13[34] ), .C(
        \R_DATA_TEMPR14[34] ), .D(\R_DATA_TEMPR15[34] ), .Y(OR4_17_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C19 (.A_DOUT({
        nc13908, nc13909, nc13910, nc13911, nc13912, nc13913, nc13914, 
        nc13915, nc13916, nc13917, nc13918, nc13919, nc13920, nc13921, 
        nc13922, nc13923, nc13924, nc13925, \R_DATA_TEMPR10[39] , 
        \R_DATA_TEMPR10[38] }), .B_DOUT({nc13926, nc13927, nc13928, 
        nc13929, nc13930, nc13931, nc13932, nc13933, nc13934, nc13935, 
        nc13936, nc13937, nc13938, nc13939, nc13940, nc13941, nc13942, 
        nc13943, nc13944, nc13945}), .DB_DETECT(\DB_DETECT[10][19] ), 
        .SB_CORRECT(\SB_CORRECT[10][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C9 (.A_DOUT({
        nc13946, nc13947, nc13948, nc13949, nc13950, nc13951, nc13952, 
        nc13953, nc13954, nc13955, nc13956, nc13957, nc13958, nc13959, 
        nc13960, nc13961, nc13962, nc13963, \R_DATA_TEMPR16[19] , 
        \R_DATA_TEMPR16[18] }), .B_DOUT({nc13964, nc13965, nc13966, 
        nc13967, nc13968, nc13969, nc13970, nc13971, nc13972, nc13973, 
        nc13974, nc13975, nc13976, nc13977, nc13978, nc13979, nc13980, 
        nc13981, nc13982, nc13983}), .DB_DETECT(\DB_DETECT[16][9] ), 
        .SB_CORRECT(\SB_CORRECT[16][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C7 (.A_DOUT({
        nc13984, nc13985, nc13986, nc13987, nc13988, nc13989, nc13990, 
        nc13991, nc13992, nc13993, nc13994, nc13995, nc13996, nc13997, 
        nc13998, nc13999, nc14000, nc14001, \R_DATA_TEMPR19[15] , 
        \R_DATA_TEMPR19[14] }), .B_DOUT({nc14002, nc14003, nc14004, 
        nc14005, nc14006, nc14007, nc14008, nc14009, nc14010, nc14011, 
        nc14012, nc14013, nc14014, nc14015, nc14016, nc14017, nc14018, 
        nc14019, nc14020, nc14021}), .DB_DETECT(\DB_DETECT[19][7] ), 
        .SB_CORRECT(\SB_CORRECT[19][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0 (.A_DOUT({
        nc14022, nc14023, nc14024, nc14025, nc14026, nc14027, nc14028, 
        nc14029, nc14030, nc14031, nc14032, nc14033, nc14034, nc14035, 
        nc14036, nc14037, nc14038, nc14039, \R_DATA_TEMPR11[1] , 
        \R_DATA_TEMPR11[0] }), .B_DOUT({nc14040, nc14041, nc14042, 
        nc14043, nc14044, nc14045, nc14046, nc14047, nc14048, nc14049, 
        nc14050, nc14051, nc14052, nc14053, nc14054, nc14055, nc14056, 
        nc14057, nc14058, nc14059}), .DB_DETECT(\DB_DETECT[11][0] ), 
        .SB_CORRECT(\SB_CORRECT[11][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C11 (.A_DOUT({
        nc14060, nc14061, nc14062, nc14063, nc14064, nc14065, nc14066, 
        nc14067, nc14068, nc14069, nc14070, nc14071, nc14072, nc14073, 
        nc14074, nc14075, nc14076, nc14077, \R_DATA_TEMPR1[23] , 
        \R_DATA_TEMPR1[22] }), .B_DOUT({nc14078, nc14079, nc14080, 
        nc14081, nc14082, nc14083, nc14084, nc14085, nc14086, nc14087, 
        nc14088, nc14089, nc14090, nc14091, nc14092, nc14093, nc14094, 
        nc14095, nc14096, nc14097}), .DB_DETECT(\DB_DETECT[1][11] ), 
        .SB_CORRECT(\SB_CORRECT[1][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C6 (.A_DOUT({nc14098, 
        nc14099, nc14100, nc14101, nc14102, nc14103, nc14104, nc14105, 
        nc14106, nc14107, nc14108, nc14109, nc14110, nc14111, nc14112, 
        nc14113, nc14114, nc14115, \R_DATA_TEMPR3[13] , 
        \R_DATA_TEMPR3[12] }), .B_DOUT({nc14116, nc14117, nc14118, 
        nc14119, nc14120, nc14121, nc14122, nc14123, nc14124, nc14125, 
        nc14126, nc14127, nc14128, nc14129, nc14130, nc14131, nc14132, 
        nc14133, nc14134, nc14135}), .DB_DETECT(\DB_DETECT[3][6] ), 
        .SB_CORRECT(\SB_CORRECT[3][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C4 (.A_DOUT({
        nc14136, nc14137, nc14138, nc14139, nc14140, nc14141, nc14142, 
        nc14143, nc14144, nc14145, nc14146, nc14147, nc14148, nc14149, 
        nc14150, nc14151, nc14152, nc14153, \R_DATA_TEMPR21[9] , 
        \R_DATA_TEMPR21[8] }), .B_DOUT({nc14154, nc14155, nc14156, 
        nc14157, nc14158, nc14159, nc14160, nc14161, nc14162, nc14163, 
        nc14164, nc14165, nc14166, nc14167, nc14168, nc14169, nc14170, 
        nc14171, nc14172, nc14173}), .DB_DETECT(\DB_DETECT[21][4] ), 
        .SB_CORRECT(\SB_CORRECT[21][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[21][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C17 (.A_DOUT({
        nc14174, nc14175, nc14176, nc14177, nc14178, nc14179, nc14180, 
        nc14181, nc14182, nc14183, nc14184, nc14185, nc14186, nc14187, 
        nc14188, nc14189, nc14190, nc14191, \R_DATA_TEMPR11[35] , 
        \R_DATA_TEMPR11[34] }), .B_DOUT({nc14192, nc14193, nc14194, 
        nc14195, nc14196, nc14197, nc14198, nc14199, nc14200, nc14201, 
        nc14202, nc14203, nc14204, nc14205, nc14206, nc14207, nc14208, 
        nc14209, nc14210, nc14211}), .DB_DETECT(\DB_DETECT[11][17] ), 
        .SB_CORRECT(\SB_CORRECT[11][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C16 (.A_DOUT({
        nc14212, nc14213, nc14214, nc14215, nc14216, nc14217, nc14218, 
        nc14219, nc14220, nc14221, nc14222, nc14223, nc14224, nc14225, 
        nc14226, nc14227, nc14228, nc14229, \R_DATA_TEMPR27[33] , 
        \R_DATA_TEMPR27[32] }), .B_DOUT({nc14230, nc14231, nc14232, 
        nc14233, nc14234, nc14235, nc14236, nc14237, nc14238, nc14239, 
        nc14240, nc14241, nc14242, nc14243, nc14244, nc14245, nc14246, 
        nc14247, nc14248, nc14249}), .DB_DETECT(\DB_DETECT[27][16] ), 
        .SB_CORRECT(\SB_CORRECT[27][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C7 (.A_DOUT({nc14250, 
        nc14251, nc14252, nc14253, nc14254, nc14255, nc14256, nc14257, 
        nc14258, nc14259, nc14260, nc14261, nc14262, nc14263, nc14264, 
        nc14265, nc14266, nc14267, \R_DATA_TEMPR4[15] , 
        \R_DATA_TEMPR4[14] }), .B_DOUT({nc14268, nc14269, nc14270, 
        nc14271, nc14272, nc14273, nc14274, nc14275, nc14276, nc14277, 
        nc14278, nc14279, nc14280, nc14281, nc14282, nc14283, nc14284, 
        nc14285, nc14286, nc14287}), .DB_DETECT(\DB_DETECT[4][7] ), 
        .SB_CORRECT(\SB_CORRECT[4][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C15 (.A_DOUT({
        nc14288, nc14289, nc14290, nc14291, nc14292, nc14293, nc14294, 
        nc14295, nc14296, nc14297, nc14298, nc14299, nc14300, nc14301, 
        nc14302, nc14303, nc14304, nc14305, \R_DATA_TEMPR5[31] , 
        \R_DATA_TEMPR5[30] }), .B_DOUT({nc14306, nc14307, nc14308, 
        nc14309, nc14310, nc14311, nc14312, nc14313, nc14314, nc14315, 
        nc14316, nc14317, nc14318, nc14319, nc14320, nc14321, nc14322, 
        nc14323, nc14324, nc14325}), .DB_DETECT(\DB_DETECT[5][15] ), 
        .SB_CORRECT(\SB_CORRECT[5][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C13 (.A_DOUT({
        nc14326, nc14327, nc14328, nc14329, nc14330, nc14331, nc14332, 
        nc14333, nc14334, nc14335, nc14336, nc14337, nc14338, nc14339, 
        nc14340, nc14341, nc14342, nc14343, \R_DATA_TEMPR19[27] , 
        \R_DATA_TEMPR19[26] }), .B_DOUT({nc14344, nc14345, nc14346, 
        nc14347, nc14348, nc14349, nc14350, nc14351, nc14352, nc14353, 
        nc14354, nc14355, nc14356, nc14357, nc14358, nc14359, nc14360, 
        nc14361, nc14362, nc14363}), .DB_DETECT(\DB_DETECT[19][13] ), 
        .SB_CORRECT(\SB_CORRECT[19][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C13 (.A_DOUT({
        nc14364, nc14365, nc14366, nc14367, nc14368, nc14369, nc14370, 
        nc14371, nc14372, nc14373, nc14374, nc14375, nc14376, nc14377, 
        nc14378, nc14379, nc14380, nc14381, \R_DATA_TEMPR22[27] , 
        \R_DATA_TEMPR22[26] }), .B_DOUT({nc14382, nc14383, nc14384, 
        nc14385, nc14386, nc14387, nc14388, nc14389, nc14390, nc14391, 
        nc14392, nc14393, nc14394, nc14395, nc14396, nc14397, nc14398, 
        nc14399, nc14400, nc14401}), .DB_DETECT(\DB_DETECT[22][13] ), 
        .SB_CORRECT(\SB_CORRECT[22][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_200 (.A(\R_DATA_TEMPR12[33] ), .B(\R_DATA_TEMPR13[33] ), 
        .C(\R_DATA_TEMPR14[33] ), .D(\R_DATA_TEMPR15[33] ), .Y(
        OR4_200_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C3 (.A_DOUT({
        nc14402, nc14403, nc14404, nc14405, nc14406, nc14407, nc14408, 
        nc14409, nc14410, nc14411, nc14412, nc14413, nc14414, nc14415, 
        nc14416, nc14417, nc14418, nc14419, \R_DATA_TEMPR17[7] , 
        \R_DATA_TEMPR17[6] }), .B_DOUT({nc14420, nc14421, nc14422, 
        nc14423, nc14424, nc14425, nc14426, nc14427, nc14428, nc14429, 
        nc14430, nc14431, nc14432, nc14433, nc14434, nc14435, nc14436, 
        nc14437, nc14438, nc14439}), .DB_DETECT(\DB_DETECT[17][3] ), 
        .SB_CORRECT(\SB_CORRECT[17][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C15 (.A_DOUT({
        nc14440, nc14441, nc14442, nc14443, nc14444, nc14445, nc14446, 
        nc14447, nc14448, nc14449, nc14450, nc14451, nc14452, nc14453, 
        nc14454, nc14455, nc14456, nc14457, \R_DATA_TEMPR27[31] , 
        \R_DATA_TEMPR27[30] }), .B_DOUT({nc14458, nc14459, nc14460, 
        nc14461, nc14462, nc14463, nc14464, nc14465, nc14466, nc14467, 
        nc14468, nc14469, nc14470, nc14471, nc14472, nc14473, nc14474, 
        nc14475, nc14476, nc14477}), .DB_DETECT(\DB_DETECT[27][15] ), 
        .SB_CORRECT(\SB_CORRECT[27][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C4 (.A_DOUT({
        nc14478, nc14479, nc14480, nc14481, nc14482, nc14483, nc14484, 
        nc14485, nc14486, nc14487, nc14488, nc14489, nc14490, nc14491, 
        nc14492, nc14493, nc14494, nc14495, \R_DATA_TEMPR28[9] , 
        \R_DATA_TEMPR28[8] }), .B_DOUT({nc14496, nc14497, nc14498, 
        nc14499, nc14500, nc14501, nc14502, nc14503, nc14504, nc14505, 
        nc14506, nc14507, nc14508, nc14509, nc14510, nc14511, nc14512, 
        nc14513, nc14514, nc14515}), .DB_DETECT(\DB_DETECT[28][4] ), 
        .SB_CORRECT(\SB_CORRECT[28][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[28][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_270 (.A(\R_DATA_TEMPR8[10] ), .B(\R_DATA_TEMPR9[10] ), .C(
        \R_DATA_TEMPR10[10] ), .D(\R_DATA_TEMPR11[10] ), .Y(OR4_270_Y));
    OR4 OR4_319 (.A(\R_DATA_TEMPR8[15] ), .B(\R_DATA_TEMPR9[15] ), .C(
        \R_DATA_TEMPR10[15] ), .D(\R_DATA_TEMPR11[15] ), .Y(OR4_319_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C18 (.A_DOUT({
        nc14516, nc14517, nc14518, nc14519, nc14520, nc14521, nc14522, 
        nc14523, nc14524, nc14525, nc14526, nc14527, nc14528, nc14529, 
        nc14530, nc14531, nc14532, nc14533, \R_DATA_TEMPR16[37] , 
        \R_DATA_TEMPR16[36] }), .B_DOUT({nc14534, nc14535, nc14536, 
        nc14537, nc14538, nc14539, nc14540, nc14541, nc14542, nc14543, 
        nc14544, nc14545, nc14546, nc14547, nc14548, nc14549, nc14550, 
        nc14551, nc14552, nc14553}), .DB_DETECT(\DB_DETECT[16][18] ), 
        .SB_CORRECT(\SB_CORRECT[16][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_192 (.A(OR4_231_Y), .B(OR4_113_Y), .C(OR4_234_Y), .D(
        OR4_104_Y), .Y(OR4_192_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C5 (.A_DOUT({nc14554, 
        nc14555, nc14556, nc14557, nc14558, nc14559, nc14560, nc14561, 
        nc14562, nc14563, nc14564, nc14565, nc14566, nc14567, nc14568, 
        nc14569, nc14570, nc14571, \R_DATA_TEMPR6[11] , 
        \R_DATA_TEMPR6[10] }), .B_DOUT({nc14572, nc14573, nc14574, 
        nc14575, nc14576, nc14577, nc14578, nc14579, nc14580, nc14581, 
        nc14582, nc14583, nc14584, nc14585, nc14586, nc14587, nc14588, 
        nc14589, nc14590, nc14591}), .DB_DETECT(\DB_DETECT[6][5] ), 
        .SB_CORRECT(\SB_CORRECT[6][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_123 (.A(\R_DATA_TEMPR12[3] ), .B(\R_DATA_TEMPR13[3] ), .C(
        \R_DATA_TEMPR14[3] ), .D(\R_DATA_TEMPR15[3] ), .Y(OR4_123_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C6 (.A_DOUT({
        nc14592, nc14593, nc14594, nc14595, nc14596, nc14597, nc14598, 
        nc14599, nc14600, nc14601, nc14602, nc14603, nc14604, nc14605, 
        nc14606, nc14607, nc14608, nc14609, \R_DATA_TEMPR25[13] , 
        \R_DATA_TEMPR25[12] }), .B_DOUT({nc14610, nc14611, nc14612, 
        nc14613, nc14614, nc14615, nc14616, nc14617, nc14618, nc14619, 
        nc14620, nc14621, nc14622, nc14623, nc14624, nc14625, nc14626, 
        nc14627, nc14628, nc14629}), .DB_DETECT(\DB_DETECT[25][6] ), 
        .SB_CORRECT(\SB_CORRECT[25][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C6 (.A_DOUT({nc14630, 
        nc14631, nc14632, nc14633, nc14634, nc14635, nc14636, nc14637, 
        nc14638, nc14639, nc14640, nc14641, nc14642, nc14643, nc14644, 
        nc14645, nc14646, nc14647, \R_DATA_TEMPR4[13] , 
        \R_DATA_TEMPR4[12] }), .B_DOUT({nc14648, nc14649, nc14650, 
        nc14651, nc14652, nc14653, nc14654, nc14655, nc14656, nc14657, 
        nc14658, nc14659, nc14660, nc14661, nc14662, nc14663, nc14664, 
        nc14665, nc14666, nc14667}), .DB_DETECT(\DB_DETECT[4][6] ), 
        .SB_CORRECT(\SB_CORRECT[4][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C17 (.A_DOUT({
        nc14668, nc14669, nc14670, nc14671, nc14672, nc14673, nc14674, 
        nc14675, nc14676, nc14677, nc14678, nc14679, nc14680, nc14681, 
        nc14682, nc14683, nc14684, nc14685, \R_DATA_TEMPR29[35] , 
        \R_DATA_TEMPR29[34] }), .B_DOUT({nc14686, nc14687, nc14688, 
        nc14689, nc14690, nc14691, nc14692, nc14693, nc14694, nc14695, 
        nc14696, nc14697, nc14698, nc14699, nc14700, nc14701, nc14702, 
        nc14703, nc14704, nc14705}), .DB_DETECT(\DB_DETECT[29][17] ), 
        .SB_CORRECT(\SB_CORRECT[29][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_206 (.A(OR4_350_Y), .B(OR4_44_Y), .C(OR4_261_Y), .D(
        OR4_215_Y), .Y(OR4_206_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C10 (.A_DOUT({
        nc14706, nc14707, nc14708, nc14709, nc14710, nc14711, nc14712, 
        nc14713, nc14714, nc14715, nc14716, nc14717, nc14718, nc14719, 
        nc14720, nc14721, nc14722, nc14723, \R_DATA_TEMPR2[21] , 
        \R_DATA_TEMPR2[20] }), .B_DOUT({nc14724, nc14725, nc14726, 
        nc14727, nc14728, nc14729, nc14730, nc14731, nc14732, nc14733, 
        nc14734, nc14735, nc14736, nc14737, nc14738, nc14739, nc14740, 
        nc14741, nc14742, nc14743}), .DB_DETECT(\DB_DETECT[2][10] ), 
        .SB_CORRECT(\SB_CORRECT[2][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C1 (.A_DOUT({
        nc14744, nc14745, nc14746, nc14747, nc14748, nc14749, nc14750, 
        nc14751, nc14752, nc14753, nc14754, nc14755, nc14756, nc14757, 
        nc14758, nc14759, nc14760, nc14761, \R_DATA_TEMPR20[3] , 
        \R_DATA_TEMPR20[2] }), .B_DOUT({nc14762, nc14763, nc14764, 
        nc14765, nc14766, nc14767, nc14768, nc14769, nc14770, nc14771, 
        nc14772, nc14773, nc14774, nc14775, nc14776, nc14777, nc14778, 
        nc14779, nc14780, nc14781}), .DB_DETECT(\DB_DETECT[20][1] ), 
        .SB_CORRECT(\SB_CORRECT[20][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C4 (.A_DOUT({nc14782, 
        nc14783, nc14784, nc14785, nc14786, nc14787, nc14788, nc14789, 
        nc14790, nc14791, nc14792, nc14793, nc14794, nc14795, nc14796, 
        nc14797, nc14798, nc14799, \R_DATA_TEMPR6[9] , 
        \R_DATA_TEMPR6[8] }), .B_DOUT({nc14800, nc14801, nc14802, 
        nc14803, nc14804, nc14805, nc14806, nc14807, nc14808, nc14809, 
        nc14810, nc14811, nc14812, nc14813, nc14814, nc14815, nc14816, 
        nc14817, nc14818, nc14819}), .DB_DETECT(\DB_DETECT[6][4] ), 
        .SB_CORRECT(\SB_CORRECT[6][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h2) )  CFG2_1 (.A(R_ADDR[16]), .B(R_ADDR[15]), .Y(
        CFG2_1_Y));
    OR4 OR4_70 (.A(\R_DATA_TEMPR24[31] ), .B(\R_DATA_TEMPR25[31] ), .C(
        \R_DATA_TEMPR26[31] ), .D(\R_DATA_TEMPR27[31] ), .Y(OR4_70_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C19 (.A_DOUT({
        nc14820, nc14821, nc14822, nc14823, nc14824, nc14825, nc14826, 
        nc14827, nc14828, nc14829, nc14830, nc14831, nc14832, nc14833, 
        nc14834, nc14835, nc14836, nc14837, \R_DATA_TEMPR14[39] , 
        \R_DATA_TEMPR14[38] }), .B_DOUT({nc14838, nc14839, nc14840, 
        nc14841, nc14842, nc14843, nc14844, nc14845, nc14846, nc14847, 
        nc14848, nc14849, nc14850, nc14851, nc14852, nc14853, nc14854, 
        nc14855, nc14856, nc14857}), .DB_DETECT(\DB_DETECT[14][19] ), 
        .SB_CORRECT(\SB_CORRECT[14][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_58 (.A(OR4_5_Y), .B(OR4_80_Y), .C(OR4_125_Y), .D(OR4_17_Y), 
        .Y(OR4_58_Y));
    OR4 OR4_276 (.A(\R_DATA_TEMPR4[27] ), .B(\R_DATA_TEMPR5[27] ), .C(
        \R_DATA_TEMPR6[27] ), .D(\R_DATA_TEMPR7[27] ), .Y(OR4_276_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C11 (.A_DOUT({
        nc14858, nc14859, nc14860, nc14861, nc14862, nc14863, nc14864, 
        nc14865, nc14866, nc14867, nc14868, nc14869, nc14870, nc14871, 
        nc14872, nc14873, nc14874, nc14875, \R_DATA_TEMPR8[23] , 
        \R_DATA_TEMPR8[22] }), .B_DOUT({nc14876, nc14877, nc14878, 
        nc14879, nc14880, nc14881, nc14882, nc14883, nc14884, nc14885, 
        nc14886, nc14887, nc14888, nc14889, nc14890, nc14891, nc14892, 
        nc14893, nc14894, nc14895}), .DB_DETECT(\DB_DETECT[8][11] ), 
        .SB_CORRECT(\SB_CORRECT[8][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_242 (.A(\R_DATA_TEMPR28[35] ), .B(\R_DATA_TEMPR29[35] ), 
        .C(\R_DATA_TEMPR30[35] ), .D(\R_DATA_TEMPR31[35] ), .Y(
        OR4_242_Y));
    OR4 OR4_77 (.A(OR4_109_Y), .B(OR4_303_Y), .C(OR4_81_Y), .D(
        OR4_250_Y), .Y(OR4_77_Y));
    OR4 OR4_299 (.A(OR4_25_Y), .B(OR2_17_Y), .C(\R_DATA_TEMPR22[34] ), 
        .D(\R_DATA_TEMPR23[34] ), .Y(OR4_299_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C19 (.A_DOUT({
        nc14896, nc14897, nc14898, nc14899, nc14900, nc14901, nc14902, 
        nc14903, nc14904, nc14905, nc14906, nc14907, nc14908, nc14909, 
        nc14910, nc14911, nc14912, nc14913, \R_DATA_TEMPR15[39] , 
        \R_DATA_TEMPR15[38] }), .B_DOUT({nc14914, nc14915, nc14916, 
        nc14917, nc14918, nc14919, nc14920, nc14921, nc14922, nc14923, 
        nc14924, nc14925, nc14926, nc14927, nc14928, nc14929, nc14930, 
        nc14931, nc14932, nc14933}), .DB_DETECT(\DB_DETECT[15][19] ), 
        .SB_CORRECT(\SB_CORRECT[15][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C6 (.A_DOUT({
        nc14934, nc14935, nc14936, nc14937, nc14938, nc14939, nc14940, 
        nc14941, nc14942, nc14943, nc14944, nc14945, nc14946, nc14947, 
        nc14948, nc14949, nc14950, nc14951, \R_DATA_TEMPR19[13] , 
        \R_DATA_TEMPR19[12] }), .B_DOUT({nc14952, nc14953, nc14954, 
        nc14955, nc14956, nc14957, nc14958, nc14959, nc14960, nc14961, 
        nc14962, nc14963, nc14964, nc14965, nc14966, nc14967, nc14968, 
        nc14969, nc14970, nc14971}), .DB_DETECT(\DB_DETECT[19][6] ), 
        .SB_CORRECT(\SB_CORRECT[19][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0 (.A_DOUT({
        nc14972, nc14973, nc14974, nc14975, nc14976, nc14977, nc14978, 
        nc14979, nc14980, nc14981, nc14982, nc14983, nc14984, nc14985, 
        nc14986, nc14987, nc14988, nc14989, \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR13[0] }), .B_DOUT({nc14990, nc14991, nc14992, 
        nc14993, nc14994, nc14995, nc14996, nc14997, nc14998, nc14999, 
        nc15000, nc15001, nc15002, nc15003, nc15004, nc15005, nc15006, 
        nc15007, nc15008, nc15009}), .DB_DETECT(\DB_DETECT[13][0] ), 
        .SB_CORRECT(\SB_CORRECT[13][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C2 (.A_DOUT({nc15010, 
        nc15011, nc15012, nc15013, nc15014, nc15015, nc15016, nc15017, 
        nc15018, nc15019, nc15020, nc15021, nc15022, nc15023, nc15024, 
        nc15025, nc15026, nc15027, \R_DATA_TEMPR0[5] , 
        \R_DATA_TEMPR0[4] }), .B_DOUT({nc15028, nc15029, nc15030, 
        nc15031, nc15032, nc15033, nc15034, nc15035, nc15036, nc15037, 
        nc15038, nc15039, nc15040, nc15041, nc15042, nc15043, nc15044, 
        nc15045, nc15046, nc15047}), .DB_DETECT(\DB_DETECT[0][2] ), 
        .SB_CORRECT(\SB_CORRECT[0][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C7 (.A_DOUT({
        nc15048, nc15049, nc15050, nc15051, nc15052, nc15053, nc15054, 
        nc15055, nc15056, nc15057, nc15058, nc15059, nc15060, nc15061, 
        nc15062, nc15063, nc15064, nc15065, \R_DATA_TEMPR10[15] , 
        \R_DATA_TEMPR10[14] }), .B_DOUT({nc15066, nc15067, nc15068, 
        nc15069, nc15070, nc15071, nc15072, nc15073, nc15074, nc15075, 
        nc15076, nc15077, nc15078, nc15079, nc15080, nc15081, nc15082, 
        nc15083, nc15084, nc15085}), .DB_DETECT(\DB_DETECT[10][7] ), 
        .SB_CORRECT(\SB_CORRECT[10][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C16 (.A_DOUT({
        nc15086, nc15087, nc15088, nc15089, nc15090, nc15091, nc15092, 
        nc15093, nc15094, nc15095, nc15096, nc15097, nc15098, nc15099, 
        nc15100, nc15101, nc15102, nc15103, \R_DATA_TEMPR22[33] , 
        \R_DATA_TEMPR22[32] }), .B_DOUT({nc15104, nc15105, nc15106, 
        nc15107, nc15108, nc15109, nc15110, nc15111, nc15112, nc15113, 
        nc15114, nc15115, nc15116, nc15117, nc15118, nc15119, nc15120, 
        nc15121, nc15122, nc15123}), .DB_DETECT(\DB_DETECT[22][16] ), 
        .SB_CORRECT(\SB_CORRECT[22][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C17 (.A_DOUT({
        nc15124, nc15125, nc15126, nc15127, nc15128, nc15129, nc15130, 
        nc15131, nc15132, nc15133, nc15134, nc15135, nc15136, nc15137, 
        nc15138, nc15139, nc15140, nc15141, \R_DATA_TEMPR31[35] , 
        \R_DATA_TEMPR31[34] }), .B_DOUT({nc15142, nc15143, nc15144, 
        nc15145, nc15146, nc15147, nc15148, nc15149, nc15150, nc15151, 
        nc15152, nc15153, nc15154, nc15155, nc15156, nc15157, nc15158, 
        nc15159, nc15160, nc15161}), .DB_DETECT(\DB_DETECT[31][17] ), 
        .SB_CORRECT(\SB_CORRECT[31][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C2 (.A_DOUT({nc15162, 
        nc15163, nc15164, nc15165, nc15166, nc15167, nc15168, nc15169, 
        nc15170, nc15171, nc15172, nc15173, nc15174, nc15175, nc15176, 
        nc15177, nc15178, nc15179, \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR4[4] }), .B_DOUT({nc15180, nc15181, nc15182, 
        nc15183, nc15184, nc15185, nc15186, nc15187, nc15188, nc15189, 
        nc15190, nc15191, nc15192, nc15193, nc15194, nc15195, nc15196, 
        nc15197, nc15198, nc15199}), .DB_DETECT(\DB_DETECT[4][2] ), 
        .SB_CORRECT(\SB_CORRECT[4][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C16 (.A_DOUT({
        nc15200, nc15201, nc15202, nc15203, nc15204, nc15205, nc15206, 
        nc15207, nc15208, nc15209, nc15210, nc15211, nc15212, nc15213, 
        nc15214, nc15215, nc15216, nc15217, \R_DATA_TEMPR4[33] , 
        \R_DATA_TEMPR4[32] }), .B_DOUT({nc15218, nc15219, nc15220, 
        nc15221, nc15222, nc15223, nc15224, nc15225, nc15226, nc15227, 
        nc15228, nc15229, nc15230, nc15231, nc15232, nc15233, nc15234, 
        nc15235, nc15236, nc15237}), .DB_DETECT(\DB_DETECT[4][16] ), 
        .SB_CORRECT(\SB_CORRECT[4][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[5]  (.A(OR4_51_Y), .B(OR4_343_Y), .C(OR4_222_Y), 
        .D(OR4_298_Y), .Y(R_DATA[5]));
    OR4 OR4_340 (.A(\R_DATA_TEMPR0[16] ), .B(\R_DATA_TEMPR1[16] ), .C(
        \R_DATA_TEMPR2[16] ), .D(\R_DATA_TEMPR3[16] ), .Y(OR4_340_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C10 (.A_DOUT({
        nc15238, nc15239, nc15240, nc15241, nc15242, nc15243, nc15244, 
        nc15245, nc15246, nc15247, nc15248, nc15249, nc15250, nc15251, 
        nc15252, nc15253, nc15254, nc15255, \R_DATA_TEMPR7[21] , 
        \R_DATA_TEMPR7[20] }), .B_DOUT({nc15256, nc15257, nc15258, 
        nc15259, nc15260, nc15261, nc15262, nc15263, nc15264, nc15265, 
        nc15266, nc15267, nc15268, nc15269, nc15270, nc15271, nc15272, 
        nc15273, nc15274, nc15275}), .DB_DETECT(\DB_DETECT[7][10] ), 
        .SB_CORRECT(\SB_CORRECT[7][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C1 (.A_DOUT({
        nc15276, nc15277, nc15278, nc15279, nc15280, nc15281, nc15282, 
        nc15283, nc15284, nc15285, nc15286, nc15287, nc15288, nc15289, 
        nc15290, nc15291, nc15292, nc15293, \R_DATA_TEMPR16[3] , 
        \R_DATA_TEMPR16[2] }), .B_DOUT({nc15294, nc15295, nc15296, 
        nc15297, nc15298, nc15299, nc15300, nc15301, nc15302, nc15303, 
        nc15304, nc15305, nc15306, nc15307, nc15308, nc15309, nc15310, 
        nc15311, nc15312, nc15313}), .DB_DETECT(\DB_DETECT[16][1] ), 
        .SB_CORRECT(\SB_CORRECT[16][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C14 (.A_DOUT({
        nc15314, nc15315, nc15316, nc15317, nc15318, nc15319, nc15320, 
        nc15321, nc15322, nc15323, nc15324, nc15325, nc15326, nc15327, 
        nc15328, nc15329, nc15330, nc15331, \R_DATA_TEMPR29[29] , 
        \R_DATA_TEMPR29[28] }), .B_DOUT({nc15332, nc15333, nc15334, 
        nc15335, nc15336, nc15337, nc15338, nc15339, nc15340, nc15341, 
        nc15342, nc15343, nc15344, nc15345, nc15346, nc15347, nc15348, 
        nc15349, nc15350, nc15351}), .DB_DETECT(\DB_DETECT[29][14] ), 
        .SB_CORRECT(\SB_CORRECT[29][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C15 (.A_DOUT({
        nc15352, nc15353, nc15354, nc15355, nc15356, nc15357, nc15358, 
        nc15359, nc15360, nc15361, nc15362, nc15363, nc15364, nc15365, 
        nc15366, nc15367, nc15368, nc15369, \R_DATA_TEMPR22[31] , 
        \R_DATA_TEMPR22[30] }), .B_DOUT({nc15370, nc15371, nc15372, 
        nc15373, nc15374, nc15375, nc15376, nc15377, nc15378, nc15379, 
        nc15380, nc15381, nc15382, nc15383, nc15384, nc15385, nc15386, 
        nc15387, nc15388, nc15389}), .DB_DETECT(\DB_DETECT[22][15] ), 
        .SB_CORRECT(\SB_CORRECT[22][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C5 (.A_DOUT({
        nc15390, nc15391, nc15392, nc15393, nc15394, nc15395, nc15396, 
        nc15397, nc15398, nc15399, nc15400, nc15401, nc15402, nc15403, 
        nc15404, nc15405, nc15406, nc15407, \R_DATA_TEMPR12[11] , 
        \R_DATA_TEMPR12[10] }), .B_DOUT({nc15408, nc15409, nc15410, 
        nc15411, nc15412, nc15413, nc15414, nc15415, nc15416, nc15417, 
        nc15418, nc15419, nc15420, nc15421, nc15422, nc15423, nc15424, 
        nc15425, nc15426, nc15427}), .DB_DETECT(\DB_DETECT[12][5] ), 
        .SB_CORRECT(\SB_CORRECT[12][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C2 (.A_DOUT({
        nc15428, nc15429, nc15430, nc15431, nc15432, nc15433, nc15434, 
        nc15435, nc15436, nc15437, nc15438, nc15439, nc15440, nc15441, 
        nc15442, nc15443, nc15444, nc15445, \R_DATA_TEMPR27[5] , 
        \R_DATA_TEMPR27[4] }), .B_DOUT({nc15446, nc15447, nc15448, 
        nc15449, nc15450, nc15451, nc15452, nc15453, nc15454, nc15455, 
        nc15456, nc15457, nc15458, nc15459, nc15460, nc15461, nc15462, 
        nc15463, nc15464, nc15465}), .DB_DETECT(\DB_DETECT[27][2] ), 
        .SB_CORRECT(\SB_CORRECT[27][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[11]  (.A(OR4_0_Y), .B(OR4_346_Y), .C(OR4_356_Y), 
        .D(OR4_237_Y), .Y(R_DATA[11]));
    OR4 OR4_122 (.A(OR4_277_Y), .B(OR2_32_Y), .C(\R_DATA_TEMPR22[39] ), 
        .D(\R_DATA_TEMPR23[39] ), .Y(OR4_122_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C7 (.A_DOUT({
        nc15466, nc15467, nc15468, nc15469, nc15470, nc15471, nc15472, 
        nc15473, nc15474, nc15475, nc15476, nc15477, nc15478, nc15479, 
        nc15480, nc15481, nc15482, nc15483, \R_DATA_TEMPR11[15] , 
        \R_DATA_TEMPR11[14] }), .B_DOUT({nc15484, nc15485, nc15486, 
        nc15487, nc15488, nc15489, nc15490, nc15491, nc15492, nc15493, 
        nc15494, nc15495, nc15496, nc15497, nc15498, nc15499, nc15500, 
        nc15501, nc15502, nc15503}), .DB_DETECT(\DB_DETECT[11][7] ), 
        .SB_CORRECT(\SB_CORRECT[11][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[9]  (.A(OR4_41_Y), .B(OR4_118_Y), .C(OR4_203_Y), 
        .D(OR4_279_Y), .Y(R_DATA[9]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C3 (.A_DOUT({
        nc15504, nc15505, nc15506, nc15507, nc15508, nc15509, nc15510, 
        nc15511, nc15512, nc15513, nc15514, nc15515, nc15516, nc15517, 
        nc15518, nc15519, nc15520, nc15521, \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR30[6] }), .B_DOUT({nc15522, nc15523, nc15524, 
        nc15525, nc15526, nc15527, nc15528, nc15529, nc15530, nc15531, 
        nc15532, nc15533, nc15534, nc15535, nc15536, nc15537, nc15538, 
        nc15539, nc15540, nc15541}), .DB_DETECT(\DB_DETECT[30][3] ), 
        .SB_CORRECT(\SB_CORRECT[30][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_18 (.A(\R_DATA_TEMPR4[35] ), .B(\R_DATA_TEMPR5[35] ), .C(
        \R_DATA_TEMPR6[35] ), .D(\R_DATA_TEMPR7[35] ), .Y(OR4_18_Y));
    OR4 OR4_34 (.A(\R_DATA_TEMPR8[35] ), .B(\R_DATA_TEMPR9[35] ), .C(
        \R_DATA_TEMPR10[35] ), .D(\R_DATA_TEMPR11[35] ), .Y(OR4_34_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C8 (.A_DOUT({
        nc15542, nc15543, nc15544, nc15545, nc15546, nc15547, nc15548, 
        nc15549, nc15550, nc15551, nc15552, nc15553, nc15554, nc15555, 
        nc15556, nc15557, nc15558, nc15559, \R_DATA_TEMPR18[17] , 
        \R_DATA_TEMPR18[16] }), .B_DOUT({nc15560, nc15561, nc15562, 
        nc15563, nc15564, nc15565, nc15566, nc15567, nc15568, nc15569, 
        nc15570, nc15571, nc15572, nc15573, nc15574, nc15575, nc15576, 
        nc15577, nc15578, nc15579}), .DB_DETECT(\DB_DETECT[18][8] ), 
        .SB_CORRECT(\SB_CORRECT[18][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1 (.A_DOUT({nc15580, 
        nc15581, nc15582, nc15583, nc15584, nc15585, nc15586, nc15587, 
        nc15588, nc15589, nc15590, nc15591, nc15592, nc15593, nc15594, 
        nc15595, nc15596, nc15597, \R_DATA_TEMPR6[3] , 
        \R_DATA_TEMPR6[2] }), .B_DOUT({nc15598, nc15599, nc15600, 
        nc15601, nc15602, nc15603, nc15604, nc15605, nc15606, nc15607, 
        nc15608, nc15609, nc15610, nc15611, nc15612, nc15613, nc15614, 
        nc15615, nc15616, nc15617}), .DB_DETECT(\DB_DETECT[6][1] ), 
        .SB_CORRECT(\SB_CORRECT[6][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C1 (.A_DOUT({
        nc15618, nc15619, nc15620, nc15621, nc15622, nc15623, nc15624, 
        nc15625, nc15626, nc15627, nc15628, nc15629, nc15630, nc15631, 
        nc15632, nc15633, nc15634, nc15635, \R_DATA_TEMPR24[3] , 
        \R_DATA_TEMPR24[2] }), .B_DOUT({nc15636, nc15637, nc15638, 
        nc15639, nc15640, nc15641, nc15642, nc15643, nc15644, nc15645, 
        nc15646, nc15647, nc15648, nc15649, nc15650, nc15651, nc15652, 
        nc15653, nc15654, nc15655}), .DB_DETECT(\DB_DETECT[24][1] ), 
        .SB_CORRECT(\SB_CORRECT[24][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C8 (.A_DOUT({
        nc15656, nc15657, nc15658, nc15659, nc15660, nc15661, nc15662, 
        nc15663, nc15664, nc15665, nc15666, nc15667, nc15668, nc15669, 
        nc15670, nc15671, nc15672, nc15673, \R_DATA_TEMPR25[17] , 
        \R_DATA_TEMPR25[16] }), .B_DOUT({nc15674, nc15675, nc15676, 
        nc15677, nc15678, nc15679, nc15680, nc15681, nc15682, nc15683, 
        nc15684, nc15685, nc15686, nc15687, nc15688, nc15689, nc15690, 
        nc15691, nc15692, nc15693}), .DB_DETECT(\DB_DETECT[25][8] ), 
        .SB_CORRECT(\SB_CORRECT[25][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C5 (.A_DOUT({
        nc15694, nc15695, nc15696, nc15697, nc15698, nc15699, nc15700, 
        nc15701, nc15702, nc15703, nc15704, nc15705, nc15706, nc15707, 
        nc15708, nc15709, nc15710, nc15711, \R_DATA_TEMPR27[11] , 
        \R_DATA_TEMPR27[10] }), .B_DOUT({nc15712, nc15713, nc15714, 
        nc15715, nc15716, nc15717, nc15718, nc15719, nc15720, nc15721, 
        nc15722, nc15723, nc15724, nc15725, nc15726, nc15727, nc15728, 
        nc15729, nc15730, nc15731}), .DB_DETECT(\DB_DETECT[27][5] ), 
        .SB_CORRECT(\SB_CORRECT[27][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C2 (.A_DOUT({
        nc15732, nc15733, nc15734, nc15735, nc15736, nc15737, nc15738, 
        nc15739, nc15740, nc15741, nc15742, nc15743, nc15744, nc15745, 
        nc15746, nc15747, nc15748, nc15749, \R_DATA_TEMPR31[5] , 
        \R_DATA_TEMPR31[4] }), .B_DOUT({nc15750, nc15751, nc15752, 
        nc15753, nc15754, nc15755, nc15756, nc15757, nc15758, nc15759, 
        nc15760, nc15761, nc15762, nc15763, nc15764, nc15765, nc15766, 
        nc15767, nc15768, nc15769}), .DB_DETECT(\DB_DETECT[31][2] ), 
        .SB_CORRECT(\SB_CORRECT[31][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[35]  (.A(OR4_27_Y), .B(OR4_204_Y), .C(OR4_352_Y), 
        .D(OR4_242_Y), .Y(R_DATA[35]));
    OR4 \OR4_R_DATA[10]  (.A(OR4_294_Y), .B(OR4_13_Y), .C(OR4_171_Y), 
        .D(OR4_33_Y), .Y(R_DATA[10]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C9 (.A_DOUT({nc15770, 
        nc15771, nc15772, nc15773, nc15774, nc15775, nc15776, nc15777, 
        nc15778, nc15779, nc15780, nc15781, nc15782, nc15783, nc15784, 
        nc15785, nc15786, nc15787, \R_DATA_TEMPR9[19] , 
        \R_DATA_TEMPR9[18] }), .B_DOUT({nc15788, nc15789, nc15790, 
        nc15791, nc15792, nc15793, nc15794, nc15795, nc15796, nc15797, 
        nc15798, nc15799, nc15800, nc15801, nc15802, nc15803, nc15804, 
        nc15805, nc15806, nc15807}), .DB_DETECT(\DB_DETECT[9][9] ), 
        .SB_CORRECT(\SB_CORRECT[9][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0 (.A_DOUT({
        nc15808, nc15809, nc15810, nc15811, nc15812, nc15813, nc15814, 
        nc15815, nc15816, nc15817, nc15818, nc15819, nc15820, nc15821, 
        nc15822, nc15823, nc15824, nc15825, \R_DATA_TEMPR19[1] , 
        \R_DATA_TEMPR19[0] }), .B_DOUT({nc15826, nc15827, nc15828, 
        nc15829, nc15830, nc15831, nc15832, nc15833, nc15834, nc15835, 
        nc15836, nc15837, nc15838, nc15839, nc15840, nc15841, nc15842, 
        nc15843, nc15844, nc15845}), .DB_DETECT(\DB_DETECT[19][0] ), 
        .SB_CORRECT(\SB_CORRECT[19][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C5 (.A_DOUT({
        nc15846, nc15847, nc15848, nc15849, nc15850, nc15851, nc15852, 
        nc15853, nc15854, nc15855, nc15856, nc15857, nc15858, nc15859, 
        nc15860, nc15861, nc15862, nc15863, \R_DATA_TEMPR25[11] , 
        \R_DATA_TEMPR25[10] }), .B_DOUT({nc15864, nc15865, nc15866, 
        nc15867, nc15868, nc15869, nc15870, nc15871, nc15872, nc15873, 
        nc15874, nc15875, nc15876, nc15877, nc15878, nc15879, nc15880, 
        nc15881, nc15882, nc15883}), .DB_DETECT(\DB_DETECT[25][5] ), 
        .SB_CORRECT(\SB_CORRECT[25][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C9 (.A_DOUT({nc15884, 
        nc15885, nc15886, nc15887, nc15888, nc15889, nc15890, nc15891, 
        nc15892, nc15893, nc15894, nc15895, nc15896, nc15897, nc15898, 
        nc15899, nc15900, nc15901, \R_DATA_TEMPR2[19] , 
        \R_DATA_TEMPR2[18] }), .B_DOUT({nc15902, nc15903, nc15904, 
        nc15905, nc15906, nc15907, nc15908, nc15909, nc15910, nc15911, 
        nc15912, nc15913, nc15914, nc15915, nc15916, nc15917, nc15918, 
        nc15919, nc15920, nc15921}), .DB_DETECT(\DB_DETECT[2][9] ), 
        .SB_CORRECT(\SB_CORRECT[2][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[1]  (.A(CFG2_2_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[1] ));
    OR4 OR4_229 (.A(\R_DATA_TEMPR4[16] ), .B(\R_DATA_TEMPR5[16] ), .C(
        \R_DATA_TEMPR6[16] ), .D(\R_DATA_TEMPR7[16] ), .Y(OR4_229_Y));
    OR4 OR4_356 (.A(\R_DATA_TEMPR24[11] ), .B(\R_DATA_TEMPR25[11] ), 
        .C(\R_DATA_TEMPR26[11] ), .D(\R_DATA_TEMPR27[11] ), .Y(
        OR4_356_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C5 (.A_DOUT({nc15922, 
        nc15923, nc15924, nc15925, nc15926, nc15927, nc15928, nc15929, 
        nc15930, nc15931, nc15932, nc15933, nc15934, nc15935, nc15936, 
        nc15937, nc15938, nc15939, \R_DATA_TEMPR0[11] , 
        \R_DATA_TEMPR0[10] }), .B_DOUT({nc15940, nc15941, nc15942, 
        nc15943, nc15944, nc15945, nc15946, nc15947, nc15948, nc15949, 
        nc15950, nc15951, nc15952, nc15953, nc15954, nc15955, nc15956, 
        nc15957, nc15958, nc15959}), .DB_DETECT(\DB_DETECT[0][5] ), 
        .SB_CORRECT(\SB_CORRECT[0][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C1 (.A_DOUT({
        nc15960, nc15961, nc15962, nc15963, nc15964, nc15965, nc15966, 
        nc15967, nc15968, nc15969, nc15970, nc15971, nc15972, nc15973, 
        nc15974, nc15975, nc15976, nc15977, \R_DATA_TEMPR25[3] , 
        \R_DATA_TEMPR25[2] }), .B_DOUT({nc15978, nc15979, nc15980, 
        nc15981, nc15982, nc15983, nc15984, nc15985, nc15986, nc15987, 
        nc15988, nc15989, nc15990, nc15991, nc15992, nc15993, nc15994, 
        nc15995, nc15996, nc15997}), .DB_DETECT(\DB_DETECT[25][1] ), 
        .SB_CORRECT(\SB_CORRECT[25][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C9 (.A_DOUT({nc15998, 
        nc15999, nc16000, nc16001, nc16002, nc16003, nc16004, nc16005, 
        nc16006, nc16007, nc16008, nc16009, nc16010, nc16011, nc16012, 
        nc16013, nc16014, nc16015, \R_DATA_TEMPR3[19] , 
        \R_DATA_TEMPR3[18] }), .B_DOUT({nc16016, nc16017, nc16018, 
        nc16019, nc16020, nc16021, nc16022, nc16023, nc16024, nc16025, 
        nc16026, nc16027, nc16028, nc16029, nc16030, nc16031, nc16032, 
        nc16033, nc16034, nc16035}), .DB_DETECT(\DB_DETECT[3][9] ), 
        .SB_CORRECT(\SB_CORRECT[3][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_261 (.A(\R_DATA_TEMPR8[7] ), .B(\R_DATA_TEMPR9[7] ), .C(
        \R_DATA_TEMPR10[7] ), .D(\R_DATA_TEMPR11[7] ), .Y(OR4_261_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C11 (.A_DOUT({
        nc16036, nc16037, nc16038, nc16039, nc16040, nc16041, nc16042, 
        nc16043, nc16044, nc16045, nc16046, nc16047, nc16048, nc16049, 
        nc16050, nc16051, nc16052, nc16053, \R_DATA_TEMPR13[23] , 
        \R_DATA_TEMPR13[22] }), .B_DOUT({nc16054, nc16055, nc16056, 
        nc16057, nc16058, nc16059, nc16060, nc16061, nc16062, nc16063, 
        nc16064, nc16065, nc16066, nc16067, nc16068, nc16069, nc16070, 
        nc16071, nc16072, nc16073}), .DB_DETECT(\DB_DETECT[13][11] ), 
        .SB_CORRECT(\SB_CORRECT[13][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C10 (.A_DOUT({
        nc16074, nc16075, nc16076, nc16077, nc16078, nc16079, nc16080, 
        nc16081, nc16082, nc16083, nc16084, nc16085, nc16086, nc16087, 
        nc16088, nc16089, nc16090, nc16091, \R_DATA_TEMPR5[21] , 
        \R_DATA_TEMPR5[20] }), .B_DOUT({nc16092, nc16093, nc16094, 
        nc16095, nc16096, nc16097, nc16098, nc16099, nc16100, nc16101, 
        nc16102, nc16103, nc16104, nc16105, nc16106, nc16107, nc16108, 
        nc16109, nc16110, nc16111}), .DB_DETECT(\DB_DETECT[5][10] ), 
        .SB_CORRECT(\SB_CORRECT[5][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_23 (.A(\R_DATA_TEMPR20[2] ), .B(\R_DATA_TEMPR21[2] ), .Y(
        OR2_23_Y));
    OR4 OR4_29 (.A(\R_DATA_TEMPR28[12] ), .B(\R_DATA_TEMPR29[12] ), .C(
        \R_DATA_TEMPR30[12] ), .D(\R_DATA_TEMPR31[12] ), .Y(OR4_29_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C8 (.A_DOUT({nc16112, 
        nc16113, nc16114, nc16115, nc16116, nc16117, nc16118, nc16119, 
        nc16120, nc16121, nc16122, nc16123, nc16124, nc16125, nc16126, 
        nc16127, nc16128, nc16129, \R_DATA_TEMPR0[17] , 
        \R_DATA_TEMPR0[16] }), .B_DOUT({nc16130, nc16131, nc16132, 
        nc16133, nc16134, nc16135, nc16136, nc16137, nc16138, nc16139, 
        nc16140, nc16141, nc16142, nc16143, nc16144, nc16145, nc16146, 
        nc16147, nc16148, nc16149}), .DB_DETECT(\DB_DETECT[0][8] ), 
        .SB_CORRECT(\SB_CORRECT[0][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[16]  (.A(OR4_160_Y), .B(OR4_2_Y), .C(OR4_63_Y), .D(
        OR4_86_Y), .Y(R_DATA[16]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C12 (.A_DOUT({
        nc16150, nc16151, nc16152, nc16153, nc16154, nc16155, nc16156, 
        nc16157, nc16158, nc16159, nc16160, nc16161, nc16162, nc16163, 
        nc16164, nc16165, nc16166, nc16167, \R_DATA_TEMPR11[25] , 
        \R_DATA_TEMPR11[24] }), .B_DOUT({nc16168, nc16169, nc16170, 
        nc16171, nc16172, nc16173, nc16174, nc16175, nc16176, nc16177, 
        nc16178, nc16179, nc16180, nc16181, nc16182, nc16183, nc16184, 
        nc16185, nc16186, nc16187}), .DB_DETECT(\DB_DETECT[11][12] ), 
        .SB_CORRECT(\SB_CORRECT[11][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C11 (.A_DOUT({
        nc16188, nc16189, nc16190, nc16191, nc16192, nc16193, nc16194, 
        nc16195, nc16196, nc16197, nc16198, nc16199, nc16200, nc16201, 
        nc16202, nc16203, nc16204, nc16205, \R_DATA_TEMPR21[23] , 
        \R_DATA_TEMPR21[22] }), .B_DOUT({nc16206, nc16207, nc16208, 
        nc16209, nc16210, nc16211, nc16212, nc16213, nc16214, nc16215, 
        nc16216, nc16217, nc16218, nc16219, nc16220, nc16221, nc16222, 
        nc16223, nc16224, nc16225}), .DB_DETECT(\DB_DETECT[21][11] ), 
        .SB_CORRECT(\SB_CORRECT[21][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[21][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C17 (.A_DOUT({
        nc16226, nc16227, nc16228, nc16229, nc16230, nc16231, nc16232, 
        nc16233, nc16234, nc16235, nc16236, nc16237, nc16238, nc16239, 
        nc16240, nc16241, nc16242, nc16243, \R_DATA_TEMPR6[35] , 
        \R_DATA_TEMPR6[34] }), .B_DOUT({nc16244, nc16245, nc16246, 
        nc16247, nc16248, nc16249, nc16250, nc16251, nc16252, nc16253, 
        nc16254, nc16255, nc16256, nc16257, nc16258, nc16259, nc16260, 
        nc16261, nc16262, nc16263}), .DB_DETECT(\DB_DETECT[6][17] ), 
        .SB_CORRECT(\SB_CORRECT[6][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_280 (.A(\R_DATA_TEMPR28[29] ), .B(\R_DATA_TEMPR29[29] ), 
        .C(\R_DATA_TEMPR30[29] ), .D(\R_DATA_TEMPR31[29] ), .Y(
        OR4_280_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C7 (.A_DOUT({nc16264, 
        nc16265, nc16266, nc16267, nc16268, nc16269, nc16270, nc16271, 
        nc16272, nc16273, nc16274, nc16275, nc16276, nc16277, nc16278, 
        nc16279, nc16280, nc16281, \R_DATA_TEMPR1[15] , 
        \R_DATA_TEMPR1[14] }), .B_DOUT({nc16282, nc16283, nc16284, 
        nc16285, nc16286, nc16287, nc16288, nc16289, nc16290, nc16291, 
        nc16292, nc16293, nc16294, nc16295, nc16296, nc16297, nc16298, 
        nc16299, nc16300, nc16301}), .DB_DETECT(\DB_DETECT[1][7] ), 
        .SB_CORRECT(\SB_CORRECT[1][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_233 (.A(\R_DATA_TEMPR4[23] ), .B(\R_DATA_TEMPR5[23] ), .C(
        \R_DATA_TEMPR6[23] ), .D(\R_DATA_TEMPR7[23] ), .Y(OR4_233_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C11 (.A_DOUT({
        nc16302, nc16303, nc16304, nc16305, nc16306, nc16307, nc16308, 
        nc16309, nc16310, nc16311, nc16312, nc16313, nc16314, nc16315, 
        nc16316, nc16317, nc16318, nc16319, \R_DATA_TEMPR31[23] , 
        \R_DATA_TEMPR31[22] }), .B_DOUT({nc16320, nc16321, nc16322, 
        nc16323, nc16324, nc16325, nc16326, nc16327, nc16328, nc16329, 
        nc16330, nc16331, nc16332, nc16333, nc16334, nc16335, nc16336, 
        nc16337, nc16338, nc16339}), .DB_DETECT(\DB_DETECT[31][11] ), 
        .SB_CORRECT(\SB_CORRECT[31][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C9 (.A_DOUT({
        nc16340, nc16341, nc16342, nc16343, nc16344, nc16345, nc16346, 
        nc16347, nc16348, nc16349, nc16350, nc16351, nc16352, nc16353, 
        nc16354, nc16355, nc16356, nc16357, \R_DATA_TEMPR31[19] , 
        \R_DATA_TEMPR31[18] }), .B_DOUT({nc16358, nc16359, nc16360, 
        nc16361, nc16362, nc16363, nc16364, nc16365, nc16366, nc16367, 
        nc16368, nc16369, nc16370, nc16371, nc16372, nc16373, nc16374, 
        nc16375, nc16376, nc16377}), .DB_DETECT(\DB_DETECT[31][9] ), 
        .SB_CORRECT(\SB_CORRECT[31][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C18 (.A_DOUT({
        nc16378, nc16379, nc16380, nc16381, nc16382, nc16383, nc16384, 
        nc16385, nc16386, nc16387, nc16388, nc16389, nc16390, nc16391, 
        nc16392, nc16393, nc16394, nc16395, \R_DATA_TEMPR17[37] , 
        \R_DATA_TEMPR17[36] }), .B_DOUT({nc16396, nc16397, nc16398, 
        nc16399, nc16400, nc16401, nc16402, nc16403, nc16404, nc16405, 
        nc16406, nc16407, nc16408, nc16409, nc16410, nc16411, nc16412, 
        nc16413, nc16414, nc16415}), .DB_DETECT(\DB_DETECT[17][18] ), 
        .SB_CORRECT(\SB_CORRECT[17][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C6 (.A_DOUT({
        nc16416, nc16417, nc16418, nc16419, nc16420, nc16421, nc16422, 
        nc16423, nc16424, nc16425, nc16426, nc16427, nc16428, nc16429, 
        nc16430, nc16431, nc16432, nc16433, \R_DATA_TEMPR26[13] , 
        \R_DATA_TEMPR26[12] }), .B_DOUT({nc16434, nc16435, nc16436, 
        nc16437, nc16438, nc16439, nc16440, nc16441, nc16442, nc16443, 
        nc16444, nc16445, nc16446, nc16447, nc16448, nc16449, nc16450, 
        nc16451, nc16452, nc16453}), .DB_DETECT(\DB_DETECT[26][6] ), 
        .SB_CORRECT(\SB_CORRECT[26][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C4 (.A_DOUT({nc16454, 
        nc16455, nc16456, nc16457, nc16458, nc16459, nc16460, nc16461, 
        nc16462, nc16463, nc16464, nc16465, nc16466, nc16467, nc16468, 
        nc16469, nc16470, nc16471, \R_DATA_TEMPR9[9] , 
        \R_DATA_TEMPR9[8] }), .B_DOUT({nc16472, nc16473, nc16474, 
        nc16475, nc16476, nc16477, nc16478, nc16479, nc16480, nc16481, 
        nc16482, nc16483, nc16484, nc16485, nc16486, nc16487, nc16488, 
        nc16489, nc16490, nc16491}), .DB_DETECT(\DB_DETECT[9][4] ), 
        .SB_CORRECT(\SB_CORRECT[9][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C7 (.A_DOUT({nc16492, 
        nc16493, nc16494, nc16495, nc16496, nc16497, nc16498, nc16499, 
        nc16500, nc16501, nc16502, nc16503, nc16504, nc16505, nc16506, 
        nc16507, nc16508, nc16509, \R_DATA_TEMPR9[15] , 
        \R_DATA_TEMPR9[14] }), .B_DOUT({nc16510, nc16511, nc16512, 
        nc16513, nc16514, nc16515, nc16516, nc16517, nc16518, nc16519, 
        nc16520, nc16521, nc16522, nc16523, nc16524, nc16525, nc16526, 
        nc16527, nc16528, nc16529}), .DB_DETECT(\DB_DETECT[9][7] ), 
        .SB_CORRECT(\SB_CORRECT[9][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C2 (.A_DOUT({
        nc16530, nc16531, nc16532, nc16533, nc16534, nc16535, nc16536, 
        nc16537, nc16538, nc16539, nc16540, nc16541, nc16542, nc16543, 
        nc16544, nc16545, nc16546, nc16547, \R_DATA_TEMPR25[5] , 
        \R_DATA_TEMPR25[4] }), .B_DOUT({nc16548, nc16549, nc16550, 
        nc16551, nc16552, nc16553, nc16554, nc16555, nc16556, nc16557, 
        nc16558, nc16559, nc16560, nc16561, nc16562, nc16563, nc16564, 
        nc16565, nc16566, nc16567}), .DB_DETECT(\DB_DETECT[25][2] ), 
        .SB_CORRECT(\SB_CORRECT[25][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C8 (.A_DOUT({nc16568, 
        nc16569, nc16570, nc16571, nc16572, nc16573, nc16574, nc16575, 
        nc16576, nc16577, nc16578, nc16579, nc16580, nc16581, nc16582, 
        nc16583, nc16584, nc16585, \R_DATA_TEMPR2[17] , 
        \R_DATA_TEMPR2[16] }), .B_DOUT({nc16586, nc16587, nc16588, 
        nc16589, nc16590, nc16591, nc16592, nc16593, nc16594, nc16595, 
        nc16596, nc16597, nc16598, nc16599, nc16600, nc16601, nc16602, 
        nc16603, nc16604, nc16605}), .DB_DETECT(\DB_DETECT[2][8] ), 
        .SB_CORRECT(\SB_CORRECT[2][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C18 (.A_DOUT({
        nc16606, nc16607, nc16608, nc16609, nc16610, nc16611, nc16612, 
        nc16613, nc16614, nc16615, nc16616, nc16617, nc16618, nc16619, 
        nc16620, nc16621, nc16622, nc16623, \R_DATA_TEMPR31[37] , 
        \R_DATA_TEMPR31[36] }), .B_DOUT({nc16624, nc16625, nc16626, 
        nc16627, nc16628, nc16629, nc16630, nc16631, nc16632, nc16633, 
        nc16634, nc16635, nc16636, nc16637, nc16638, nc16639, nc16640, 
        nc16641, nc16642, nc16643}), .DB_DETECT(\DB_DETECT[31][18] ), 
        .SB_CORRECT(\SB_CORRECT[31][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C15 (.A_DOUT({
        nc16644, nc16645, nc16646, nc16647, nc16648, nc16649, nc16650, 
        nc16651, nc16652, nc16653, nc16654, nc16655, nc16656, nc16657, 
        nc16658, nc16659, nc16660, nc16661, \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR1[30] }), .B_DOUT({nc16662, nc16663, nc16664, 
        nc16665, nc16666, nc16667, nc16668, nc16669, nc16670, nc16671, 
        nc16672, nc16673, nc16674, nc16675, nc16676, nc16677, nc16678, 
        nc16679, nc16680, nc16681}), .DB_DETECT(\DB_DETECT[1][15] ), 
        .SB_CORRECT(\SB_CORRECT[1][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_286 (.A(\R_DATA_TEMPR0[14] ), .B(\R_DATA_TEMPR1[14] ), .C(
        \R_DATA_TEMPR2[14] ), .D(\R_DATA_TEMPR3[14] ), .Y(OR4_286_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C6 (.A_DOUT({
        nc16682, nc16683, nc16684, nc16685, nc16686, nc16687, nc16688, 
        nc16689, nc16690, nc16691, nc16692, nc16693, nc16694, nc16695, 
        nc16696, nc16697, nc16698, nc16699, \R_DATA_TEMPR18[13] , 
        \R_DATA_TEMPR18[12] }), .B_DOUT({nc16700, nc16701, nc16702, 
        nc16703, nc16704, nc16705, nc16706, nc16707, nc16708, nc16709, 
        nc16710, nc16711, nc16712, nc16713, nc16714, nc16715, nc16716, 
        nc16717, nc16718, nc16719}), .DB_DETECT(\DB_DETECT[18][6] ), 
        .SB_CORRECT(\SB_CORRECT[18][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_78 (.A(\R_DATA_TEMPR12[9] ), .B(\R_DATA_TEMPR13[9] ), .C(
        \R_DATA_TEMPR14[9] ), .D(\R_DATA_TEMPR15[9] ), .Y(OR4_78_Y));
    OR4 \OR4_R_DATA[8]  (.A(OR4_174_Y), .B(OR4_214_Y), .C(OR4_134_Y), 
        .D(OR4_269_Y), .Y(R_DATA[8]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C13 (.A_DOUT({
        nc16720, nc16721, nc16722, nc16723, nc16724, nc16725, nc16726, 
        nc16727, nc16728, nc16729, nc16730, nc16731, nc16732, nc16733, 
        nc16734, nc16735, nc16736, nc16737, \R_DATA_TEMPR29[27] , 
        \R_DATA_TEMPR29[26] }), .B_DOUT({nc16738, nc16739, nc16740, 
        nc16741, nc16742, nc16743, nc16744, nc16745, nc16746, nc16747, 
        nc16748, nc16749, nc16750, nc16751, nc16752, nc16753, nc16754, 
        nc16755, nc16756, nc16757}), .DB_DETECT(\DB_DETECT[29][13] ), 
        .SB_CORRECT(\SB_CORRECT[29][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_154 (.A(\R_DATA_TEMPR4[20] ), .B(\R_DATA_TEMPR5[20] ), .C(
        \R_DATA_TEMPR6[20] ), .D(\R_DATA_TEMPR7[20] ), .Y(OR4_154_Y));
    OR2 OR2_21 (.A(\R_DATA_TEMPR20[8] ), .B(\R_DATA_TEMPR21[8] ), .Y(
        OR2_21_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C13 (.A_DOUT({
        nc16758, nc16759, nc16760, nc16761, nc16762, nc16763, nc16764, 
        nc16765, nc16766, nc16767, nc16768, nc16769, nc16770, nc16771, 
        nc16772, nc16773, nc16774, nc16775, \R_DATA_TEMPR30[27] , 
        \R_DATA_TEMPR30[26] }), .B_DOUT({nc16776, nc16777, nc16778, 
        nc16779, nc16780, nc16781, nc16782, nc16783, nc16784, nc16785, 
        nc16786, nc16787, nc16788, nc16789, nc16790, nc16791, nc16792, 
        nc16793, nc16794, nc16795}), .DB_DETECT(\DB_DETECT[30][13] ), 
        .SB_CORRECT(\SB_CORRECT[30][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_22 (.A(\R_DATA_TEMPR28[39] ), .B(\R_DATA_TEMPR29[39] ), .C(
        \R_DATA_TEMPR30[39] ), .D(\R_DATA_TEMPR31[39] ), .Y(OR4_22_Y));
    OR4 OR4_143 (.A(\R_DATA_TEMPR28[28] ), .B(\R_DATA_TEMPR29[28] ), 
        .C(\R_DATA_TEMPR30[28] ), .D(\R_DATA_TEMPR31[28] ), .Y(
        OR4_143_Y));
    OR4 OR4_213 (.A(OR4_62_Y), .B(OR2_16_Y), .C(\R_DATA_TEMPR22[22] ), 
        .D(\R_DATA_TEMPR23[22] ), .Y(OR4_213_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C1 (.A_DOUT({
        nc16796, nc16797, nc16798, nc16799, nc16800, nc16801, nc16802, 
        nc16803, nc16804, nc16805, nc16806, nc16807, nc16808, nc16809, 
        nc16810, nc16811, nc16812, nc16813, \R_DATA_TEMPR17[3] , 
        \R_DATA_TEMPR17[2] }), .B_DOUT({nc16814, nc16815, nc16816, 
        nc16817, nc16818, nc16819, nc16820, nc16821, nc16822, nc16823, 
        nc16824, nc16825, nc16826, nc16827, nc16828, nc16829, nc16830, 
        nc16831, nc16832, nc16833}), .DB_DETECT(\DB_DETECT[17][1] ), 
        .SB_CORRECT(\SB_CORRECT[17][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0 (.A_DOUT({
        nc16834, nc16835, nc16836, nc16837, nc16838, nc16839, nc16840, 
        nc16841, nc16842, nc16843, nc16844, nc16845, nc16846, nc16847, 
        nc16848, nc16849, nc16850, nc16851, \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR10[0] }), .B_DOUT({nc16852, nc16853, nc16854, 
        nc16855, nc16856, nc16857, nc16858, nc16859, nc16860, nc16861, 
        nc16862, nc16863, nc16864, nc16865, nc16866, nc16867, nc16868, 
        nc16869, nc16870, nc16871}), .DB_DETECT(\DB_DETECT[10][0] ), 
        .SB_CORRECT(\SB_CORRECT[10][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C8 (.A_DOUT({
        nc16872, nc16873, nc16874, nc16875, nc16876, nc16877, nc16878, 
        nc16879, nc16880, nc16881, nc16882, nc16883, nc16884, nc16885, 
        nc16886, nc16887, nc16888, nc16889, \R_DATA_TEMPR31[17] , 
        \R_DATA_TEMPR31[16] }), .B_DOUT({nc16890, nc16891, nc16892, 
        nc16893, nc16894, nc16895, nc16896, nc16897, nc16898, nc16899, 
        nc16900, nc16901, nc16902, nc16903, nc16904, nc16905, nc16906, 
        nc16907, nc16908, nc16909}), .DB_DETECT(\DB_DETECT[31][8] ), 
        .SB_CORRECT(\SB_CORRECT[31][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C8 (.A_DOUT({nc16910, 
        nc16911, nc16912, nc16913, nc16914, nc16915, nc16916, nc16917, 
        nc16918, nc16919, nc16920, nc16921, nc16922, nc16923, nc16924, 
        nc16925, nc16926, nc16927, \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR1[16] }), .B_DOUT({nc16928, nc16929, nc16930, 
        nc16931, nc16932, nc16933, nc16934, nc16935, nc16936, nc16937, 
        nc16938, nc16939, nc16940, nc16941, nc16942, nc16943, nc16944, 
        nc16945, nc16946, nc16947}), .DB_DETECT(\DB_DETECT[1][8] ), 
        .SB_CORRECT(\SB_CORRECT[1][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_201 (.A(\R_DATA_TEMPR0[31] ), .B(\R_DATA_TEMPR1[31] ), .C(
        \R_DATA_TEMPR2[31] ), .D(\R_DATA_TEMPR3[31] ), .Y(OR4_201_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C7 (.A_DOUT({nc16948, 
        nc16949, nc16950, nc16951, nc16952, nc16953, nc16954, nc16955, 
        nc16956, nc16957, nc16958, nc16959, nc16960, nc16961, nc16962, 
        nc16963, nc16964, nc16965, \R_DATA_TEMPR7[15] , 
        \R_DATA_TEMPR7[14] }), .B_DOUT({nc16966, nc16967, nc16968, 
        nc16969, nc16970, nc16971, nc16972, nc16973, nc16974, nc16975, 
        nc16976, nc16977, nc16978, nc16979, nc16980, nc16981, nc16982, 
        nc16983, nc16984, nc16985}), .DB_DETECT(\DB_DETECT[7][7] ), 
        .SB_CORRECT(\SB_CORRECT[7][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_13 (.A(\R_DATA_TEMPR20[18] ), .B(\R_DATA_TEMPR21[18] ), .Y(
        OR2_13_Y));
    OR4 OR4_6 (.A(\R_DATA_TEMPR12[1] ), .B(\R_DATA_TEMPR13[1] ), .C(
        \R_DATA_TEMPR14[1] ), .D(\R_DATA_TEMPR15[1] ), .Y(OR4_6_Y));
    OR4 OR4_271 (.A(\R_DATA_TEMPR28[34] ), .B(\R_DATA_TEMPR29[34] ), 
        .C(\R_DATA_TEMPR30[34] ), .D(\R_DATA_TEMPR31[34] ), .Y(
        OR4_271_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C8 (.A_DOUT({nc16986, 
        nc16987, nc16988, nc16989, nc16990, nc16991, nc16992, nc16993, 
        nc16994, nc16995, nc16996, nc16997, nc16998, nc16999, nc17000, 
        nc17001, nc17002, nc17003, \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR4[16] }), .B_DOUT({nc17004, nc17005, nc17006, 
        nc17007, nc17008, nc17009, nc17010, nc17011, nc17012, nc17013, 
        nc17014, nc17015, nc17016, nc17017, nc17018, nc17019, nc17020, 
        nc17021, nc17022, nc17023}), .DB_DETECT(\DB_DETECT[4][8] ), 
        .SB_CORRECT(\SB_CORRECT[4][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C10 (.A_DOUT({
        nc17024, nc17025, nc17026, nc17027, nc17028, nc17029, nc17030, 
        nc17031, nc17032, nc17033, nc17034, nc17035, nc17036, nc17037, 
        nc17038, nc17039, nc17040, nc17041, \R_DATA_TEMPR16[21] , 
        \R_DATA_TEMPR16[20] }), .B_DOUT({nc17042, nc17043, nc17044, 
        nc17045, nc17046, nc17047, nc17048, nc17049, nc17050, nc17051, 
        nc17052, nc17053, nc17054, nc17055, nc17056, nc17057, nc17058, 
        nc17059, nc17060, nc17061}), .DB_DETECT(\DB_DETECT[16][10] ), 
        .SB_CORRECT(\SB_CORRECT[16][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0 (.A_DOUT({
        nc17062, nc17063, nc17064, nc17065, nc17066, nc17067, nc17068, 
        nc17069, nc17070, nc17071, nc17072, nc17073, nc17074, nc17075, 
        nc17076, nc17077, nc17078, nc17079, \R_DATA_TEMPR26[1] , 
        \R_DATA_TEMPR26[0] }), .B_DOUT({nc17080, nc17081, nc17082, 
        nc17083, nc17084, nc17085, nc17086, nc17087, nc17088, nc17089, 
        nc17090, nc17091, nc17092, nc17093, nc17094, nc17095, nc17096, 
        nc17097, nc17098, nc17099}), .DB_DETECT(\DB_DETECT[26][0] ), 
        .SB_CORRECT(\SB_CORRECT[26][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C18 (.A_DOUT({
        nc17100, nc17101, nc17102, nc17103, nc17104, nc17105, nc17106, 
        nc17107, nc17108, nc17109, nc17110, nc17111, nc17112, nc17113, 
        nc17114, nc17115, nc17116, nc17117, \R_DATA_TEMPR12[37] , 
        \R_DATA_TEMPR12[36] }), .B_DOUT({nc17118, nc17119, nc17120, 
        nc17121, nc17122, nc17123, nc17124, nc17125, nc17126, nc17127, 
        nc17128, nc17129, nc17130, nc17131, nc17132, nc17133, nc17134, 
        nc17135, nc17136, nc17137}), .DB_DETECT(\DB_DETECT[12][18] ), 
        .SB_CORRECT(\SB_CORRECT[12][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C9 (.A_DOUT({
        nc17138, nc17139, nc17140, nc17141, nc17142, nc17143, nc17144, 
        nc17145, nc17146, nc17147, nc17148, nc17149, nc17150, nc17151, 
        nc17152, nc17153, nc17154, nc17155, \R_DATA_TEMPR17[19] , 
        \R_DATA_TEMPR17[18] }), .B_DOUT({nc17156, nc17157, nc17158, 
        nc17159, nc17160, nc17161, nc17162, nc17163, nc17164, nc17165, 
        nc17166, nc17167, nc17168, nc17169, nc17170, nc17171, nc17172, 
        nc17173, nc17174, nc17175}), .DB_DETECT(\DB_DETECT[17][9] ), 
        .SB_CORRECT(\SB_CORRECT[17][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C4 (.A_DOUT({
        nc17176, nc17177, nc17178, nc17179, nc17180, nc17181, nc17182, 
        nc17183, nc17184, nc17185, nc17186, nc17187, nc17188, nc17189, 
        nc17190, nc17191, nc17192, nc17193, \R_DATA_TEMPR13[9] , 
        \R_DATA_TEMPR13[8] }), .B_DOUT({nc17194, nc17195, nc17196, 
        nc17197, nc17198, nc17199, nc17200, nc17201, nc17202, nc17203, 
        nc17204, nc17205, nc17206, nc17207, nc17208, nc17209, nc17210, 
        nc17211, nc17212, nc17213}), .DB_DETECT(\DB_DETECT[13][4] ), 
        .SB_CORRECT(\SB_CORRECT[13][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C15 (.A_DOUT({
        nc17214, nc17215, nc17216, nc17217, nc17218, nc17219, nc17220, 
        nc17221, nc17222, nc17223, nc17224, nc17225, nc17226, nc17227, 
        nc17228, nc17229, nc17230, nc17231, \R_DATA_TEMPR16[31] , 
        \R_DATA_TEMPR16[30] }), .B_DOUT({nc17232, nc17233, nc17234, 
        nc17235, nc17236, nc17237, nc17238, nc17239, nc17240, nc17241, 
        nc17242, nc17243, nc17244, nc17245, nc17246, nc17247, nc17248, 
        nc17249, nc17250, nc17251}), .DB_DETECT(\DB_DETECT[16][15] ), 
        .SB_CORRECT(\SB_CORRECT[16][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C11 (.A_DOUT({
        nc17252, nc17253, nc17254, nc17255, nc17256, nc17257, nc17258, 
        nc17259, nc17260, nc17261, nc17262, nc17263, nc17264, nc17265, 
        nc17266, nc17267, nc17268, nc17269, \R_DATA_TEMPR10[23] , 
        \R_DATA_TEMPR10[22] }), .B_DOUT({nc17270, nc17271, nc17272, 
        nc17273, nc17274, nc17275, nc17276, nc17277, nc17278, nc17279, 
        nc17280, nc17281, nc17282, nc17283, nc17284, nc17285, nc17286, 
        nc17287, nc17288, nc17289}), .DB_DETECT(\DB_DETECT[10][11] ), 
        .SB_CORRECT(\SB_CORRECT[10][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C16 (.A_DOUT({
        nc17290, nc17291, nc17292, nc17293, nc17294, nc17295, nc17296, 
        nc17297, nc17298, nc17299, nc17300, nc17301, nc17302, nc17303, 
        nc17304, nc17305, nc17306, nc17307, \R_DATA_TEMPR3[33] , 
        \R_DATA_TEMPR3[32] }), .B_DOUT({nc17308, nc17309, nc17310, 
        nc17311, nc17312, nc17313, nc17314, nc17315, nc17316, nc17317, 
        nc17318, nc17319, nc17320, nc17321, nc17322, nc17323, nc17324, 
        nc17325, nc17326, nc17327}), .DB_DETECT(\DB_DETECT[3][16] ), 
        .SB_CORRECT(\SB_CORRECT[3][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C15 (.A_DOUT({
        nc17328, nc17329, nc17330, nc17331, nc17332, nc17333, nc17334, 
        nc17335, nc17336, nc17337, nc17338, nc17339, nc17340, nc17341, 
        nc17342, nc17343, nc17344, nc17345, \R_DATA_TEMPR8[31] , 
        \R_DATA_TEMPR8[30] }), .B_DOUT({nc17346, nc17347, nc17348, 
        nc17349, nc17350, nc17351, nc17352, nc17353, nc17354, nc17355, 
        nc17356, nc17357, nc17358, nc17359, nc17360, nc17361, nc17362, 
        nc17363, nc17364, nc17365}), .DB_DETECT(\DB_DETECT[8][15] ), 
        .SB_CORRECT(\SB_CORRECT[8][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C3 (.A_DOUT({
        nc17366, nc17367, nc17368, nc17369, nc17370, nc17371, nc17372, 
        nc17373, nc17374, nc17375, nc17376, nc17377, nc17378, nc17379, 
        nc17380, nc17381, nc17382, nc17383, \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR15[6] }), .B_DOUT({nc17384, nc17385, nc17386, 
        nc17387, nc17388, nc17389, nc17390, nc17391, nc17392, nc17393, 
        nc17394, nc17395, nc17396, nc17397, nc17398, nc17399, nc17400, 
        nc17401, nc17402, nc17403}), .DB_DETECT(\DB_DETECT[15][3] ), 
        .SB_CORRECT(\SB_CORRECT[15][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C4 (.A_DOUT({
        nc17404, nc17405, nc17406, nc17407, nc17408, nc17409, nc17410, 
        nc17411, nc17412, nc17413, nc17414, nc17415, nc17416, nc17417, 
        nc17418, nc17419, nc17420, nc17421, \R_DATA_TEMPR10[9] , 
        \R_DATA_TEMPR10[8] }), .B_DOUT({nc17422, nc17423, nc17424, 
        nc17425, nc17426, nc17427, nc17428, nc17429, nc17430, nc17431, 
        nc17432, nc17433, nc17434, nc17435, nc17436, nc17437, nc17438, 
        nc17439, nc17440, nc17441}), .DB_DETECT(\DB_DETECT[10][4] ), 
        .SB_CORRECT(\SB_CORRECT[10][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C16 (.A_DOUT({
        nc17442, nc17443, nc17444, nc17445, nc17446, nc17447, nc17448, 
        nc17449, nc17450, nc17451, nc17452, nc17453, nc17454, nc17455, 
        nc17456, nc17457, nc17458, nc17459, \R_DATA_TEMPR29[33] , 
        \R_DATA_TEMPR29[32] }), .B_DOUT({nc17460, nc17461, nc17462, 
        nc17463, nc17464, nc17465, nc17466, nc17467, nc17468, nc17469, 
        nc17470, nc17471, nc17472, nc17473, nc17474, nc17475, nc17476, 
        nc17477, nc17478, nc17479}), .DB_DETECT(\DB_DETECT[29][16] ), 
        .SB_CORRECT(\SB_CORRECT[29][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C9 (.A_DOUT({nc17480, 
        nc17481, nc17482, nc17483, nc17484, nc17485, nc17486, nc17487, 
        nc17488, nc17489, nc17490, nc17491, nc17492, nc17493, nc17494, 
        nc17495, nc17496, nc17497, \R_DATA_TEMPR1[19] , 
        \R_DATA_TEMPR1[18] }), .B_DOUT({nc17498, nc17499, nc17500, 
        nc17501, nc17502, nc17503, nc17504, nc17505, nc17506, nc17507, 
        nc17508, nc17509, nc17510, nc17511, nc17512, nc17513, nc17514, 
        nc17515, nc17516, nc17517}), .DB_DETECT(\DB_DETECT[1][9] ), 
        .SB_CORRECT(\SB_CORRECT[1][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[17]  (.A(OR4_77_Y), .B(OR4_244_Y), .C(OR4_339_Y), 
        .D(OR4_12_Y), .Y(R_DATA[17]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C8 (.A_DOUT({
        nc17518, nc17519, nc17520, nc17521, nc17522, nc17523, nc17524, 
        nc17525, nc17526, nc17527, nc17528, nc17529, nc17530, nc17531, 
        nc17532, nc17533, nc17534, nc17535, \R_DATA_TEMPR16[17] , 
        \R_DATA_TEMPR16[16] }), .B_DOUT({nc17536, nc17537, nc17538, 
        nc17539, nc17540, nc17541, nc17542, nc17543, nc17544, nc17545, 
        nc17546, nc17547, nc17548, nc17549, nc17550, nc17551, nc17552, 
        nc17553, nc17554, nc17555}), .DB_DETECT(\DB_DETECT[16][8] ), 
        .SB_CORRECT(\SB_CORRECT[16][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_142 (.A(\R_DATA_TEMPR24[36] ), .B(\R_DATA_TEMPR25[36] ), 
        .C(\R_DATA_TEMPR26[36] ), .D(\R_DATA_TEMPR27[36] ), .Y(
        OR4_142_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C13 (.A_DOUT({
        nc17556, nc17557, nc17558, nc17559, nc17560, nc17561, nc17562, 
        nc17563, nc17564, nc17565, nc17566, nc17567, nc17568, nc17569, 
        nc17570, nc17571, nc17572, nc17573, \R_DATA_TEMPR6[27] , 
        \R_DATA_TEMPR6[26] }), .B_DOUT({nc17574, nc17575, nc17576, 
        nc17577, nc17578, nc17579, nc17580, nc17581, nc17582, nc17583, 
        nc17584, nc17585, nc17586, nc17587, nc17588, nc17589, nc17590, 
        nc17591, nc17592, nc17593}), .DB_DETECT(\DB_DETECT[6][13] ), 
        .SB_CORRECT(\SB_CORRECT[6][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C7 (.A_DOUT({
        nc17594, nc17595, nc17596, nc17597, nc17598, nc17599, nc17600, 
        nc17601, nc17602, nc17603, nc17604, nc17605, nc17606, nc17607, 
        nc17608, nc17609, nc17610, nc17611, \R_DATA_TEMPR18[15] , 
        \R_DATA_TEMPR18[14] }), .B_DOUT({nc17612, nc17613, nc17614, 
        nc17615, nc17616, nc17617, nc17618, nc17619, nc17620, nc17621, 
        nc17622, nc17623, nc17624, nc17625, nc17626, nc17627, nc17628, 
        nc17629, nc17630, nc17631}), .DB_DETECT(\DB_DETECT[18][7] ), 
        .SB_CORRECT(\SB_CORRECT[18][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C15 (.A_DOUT({
        nc17632, nc17633, nc17634, nc17635, nc17636, nc17637, nc17638, 
        nc17639, nc17640, nc17641, nc17642, nc17643, nc17644, nc17645, 
        nc17646, nc17647, nc17648, nc17649, \R_DATA_TEMPR29[31] , 
        \R_DATA_TEMPR29[30] }), .B_DOUT({nc17650, nc17651, nc17652, 
        nc17653, nc17654, nc17655, nc17656, nc17657, nc17658, nc17659, 
        nc17660, nc17661, nc17662, nc17663, nc17664, nc17665, nc17666, 
        nc17667, nc17668, nc17669}), .DB_DETECT(\DB_DETECT[29][15] ), 
        .SB_CORRECT(\SB_CORRECT[29][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C12 (.A_DOUT({
        nc17670, nc17671, nc17672, nc17673, nc17674, nc17675, nc17676, 
        nc17677, nc17678, nc17679, nc17680, nc17681, nc17682, nc17683, 
        nc17684, nc17685, nc17686, nc17687, \R_DATA_TEMPR9[25] , 
        \R_DATA_TEMPR9[24] }), .B_DOUT({nc17688, nc17689, nc17690, 
        nc17691, nc17692, nc17693, nc17694, nc17695, nc17696, nc17697, 
        nc17698, nc17699, nc17700, nc17701, nc17702, nc17703, nc17704, 
        nc17705, nc17706, nc17707}), .DB_DETECT(\DB_DETECT[9][12] ), 
        .SB_CORRECT(\SB_CORRECT[9][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C7 (.A_DOUT({
        nc17708, nc17709, nc17710, nc17711, nc17712, nc17713, nc17714, 
        nc17715, nc17716, nc17717, nc17718, nc17719, nc17720, nc17721, 
        nc17722, nc17723, nc17724, nc17725, \R_DATA_TEMPR24[15] , 
        \R_DATA_TEMPR24[14] }), .B_DOUT({nc17726, nc17727, nc17728, 
        nc17729, nc17730, nc17731, nc17732, nc17733, nc17734, nc17735, 
        nc17736, nc17737, nc17738, nc17739, nc17740, nc17741, nc17742, 
        nc17743, nc17744, nc17745}), .DB_DETECT(\DB_DETECT[24][7] ), 
        .SB_CORRECT(\SB_CORRECT[24][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C14 (.A_DOUT({
        nc17746, nc17747, nc17748, nc17749, nc17750, nc17751, nc17752, 
        nc17753, nc17754, nc17755, nc17756, nc17757, nc17758, nc17759, 
        nc17760, nc17761, nc17762, nc17763, \R_DATA_TEMPR4[29] , 
        \R_DATA_TEMPR4[28] }), .B_DOUT({nc17764, nc17765, nc17766, 
        nc17767, nc17768, nc17769, nc17770, nc17771, nc17772, nc17773, 
        nc17774, nc17775, nc17776, nc17777, nc17778, nc17779, nc17780, 
        nc17781, nc17782, nc17783}), .DB_DETECT(\DB_DETECT[4][14] ), 
        .SB_CORRECT(\SB_CORRECT[4][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_11 (.A(\R_DATA_TEMPR20[30] ), .B(\R_DATA_TEMPR21[30] ), .Y(
        OR2_11_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C5 (.A_DOUT({
        nc17784, nc17785, nc17786, nc17787, nc17788, nc17789, nc17790, 
        nc17791, nc17792, nc17793, nc17794, nc17795, nc17796, nc17797, 
        nc17798, nc17799, nc17800, nc17801, \R_DATA_TEMPR13[11] , 
        \R_DATA_TEMPR13[10] }), .B_DOUT({nc17802, nc17803, nc17804, 
        nc17805, nc17806, nc17807, nc17808, nc17809, nc17810, nc17811, 
        nc17812, nc17813, nc17814, nc17815, nc17816, nc17817, nc17818, 
        nc17819, nc17820, nc17821}), .DB_DETECT(\DB_DETECT[13][5] ), 
        .SB_CORRECT(\SB_CORRECT[13][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1 (.A_DOUT({
        nc17822, nc17823, nc17824, nc17825, nc17826, nc17827, nc17828, 
        nc17829, nc17830, nc17831, nc17832, nc17833, nc17834, nc17835, 
        nc17836, nc17837, nc17838, nc17839, \R_DATA_TEMPR12[3] , 
        \R_DATA_TEMPR12[2] }), .B_DOUT({nc17840, nc17841, nc17842, 
        nc17843, nc17844, nc17845, nc17846, nc17847, nc17848, nc17849, 
        nc17850, nc17851, nc17852, nc17853, nc17854, nc17855, nc17856, 
        nc17857, nc17858, nc17859}), .DB_DETECT(\DB_DETECT[12][1] ), 
        .SB_CORRECT(\SB_CORRECT[12][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C19 (.A_DOUT({
        nc17860, nc17861, nc17862, nc17863, nc17864, nc17865, nc17866, 
        nc17867, nc17868, nc17869, nc17870, nc17871, nc17872, nc17873, 
        nc17874, nc17875, nc17876, nc17877, \R_DATA_TEMPR31[39] , 
        \R_DATA_TEMPR31[38] }), .B_DOUT({nc17878, nc17879, nc17880, 
        nc17881, nc17882, nc17883, nc17884, nc17885, nc17886, nc17887, 
        nc17888, nc17889, nc17890, nc17891, nc17892, nc17893, nc17894, 
        nc17895, nc17896, nc17897}), .DB_DETECT(\DB_DETECT[31][19] ), 
        .SB_CORRECT(\SB_CORRECT[31][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_55 (.A(\R_DATA_TEMPR28[6] ), .B(\R_DATA_TEMPR29[6] ), .C(
        \R_DATA_TEMPR30[6] ), .D(\R_DATA_TEMPR31[6] ), .Y(OR4_55_Y));
    OR4 OR4_301 (.A(OR4_54_Y), .B(OR4_357_Y), .C(OR4_348_Y), .D(
        OR4_200_Y), .Y(OR4_301_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C10 (.A_DOUT({
        nc17898, nc17899, nc17900, nc17901, nc17902, nc17903, nc17904, 
        nc17905, nc17906, nc17907, nc17908, nc17909, nc17910, nc17911, 
        nc17912, nc17913, nc17914, nc17915, \R_DATA_TEMPR1[21] , 
        \R_DATA_TEMPR1[20] }), .B_DOUT({nc17916, nc17917, nc17918, 
        nc17919, nc17920, nc17921, nc17922, nc17923, nc17924, nc17925, 
        nc17926, nc17927, nc17928, nc17929, nc17930, nc17931, nc17932, 
        nc17933, nc17934, nc17935}), .DB_DETECT(\DB_DETECT[1][10] ), 
        .SB_CORRECT(\SB_CORRECT[1][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_249 (.A(\R_DATA_TEMPR0[24] ), .B(\R_DATA_TEMPR1[24] ), .C(
        \R_DATA_TEMPR2[24] ), .D(\R_DATA_TEMPR3[24] ), .Y(OR4_249_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C11 (.A_DOUT({
        nc17936, nc17937, nc17938, nc17939, nc17940, nc17941, nc17942, 
        nc17943, nc17944, nc17945, nc17946, nc17947, nc17948, nc17949, 
        nc17950, nc17951, nc17952, nc17953, \R_DATA_TEMPR14[23] , 
        \R_DATA_TEMPR14[22] }), .B_DOUT({nc17954, nc17955, nc17956, 
        nc17957, nc17958, nc17959, nc17960, nc17961, nc17962, nc17963, 
        nc17964, nc17965, nc17966, nc17967, nc17968, nc17969, nc17970, 
        nc17971, nc17972, nc17973}), .DB_DETECT(\DB_DETECT[14][11] ), 
        .SB_CORRECT(\SB_CORRECT[14][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C7 (.A_DOUT({nc17974, 
        nc17975, nc17976, nc17977, nc17978, nc17979, nc17980, nc17981, 
        nc17982, nc17983, nc17984, nc17985, nc17986, nc17987, nc17988, 
        nc17989, nc17990, nc17991, \R_DATA_TEMPR3[15] , 
        \R_DATA_TEMPR3[14] }), .B_DOUT({nc17992, nc17993, nc17994, 
        nc17995, nc17996, nc17997, nc17998, nc17999, nc18000, nc18001, 
        nc18002, nc18003, nc18004, nc18005, nc18006, nc18007, nc18008, 
        nc18009, nc18010, nc18011}), .DB_DETECT(\DB_DETECT[3][7] ), 
        .SB_CORRECT(\SB_CORRECT[3][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[38]  (.A(OR4_60_Y), .B(OR4_15_Y), .C(OR4_208_Y), 
        .D(OR4_260_Y), .Y(R_DATA[38]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0 (.A_DOUT({nc18012, 
        nc18013, nc18014, nc18015, nc18016, nc18017, nc18018, nc18019, 
        nc18020, nc18021, nc18022, nc18023, nc18024, nc18025, nc18026, 
        nc18027, nc18028, nc18029, \R_DATA_TEMPR0[1] , 
        \R_DATA_TEMPR0[0] }), .B_DOUT({nc18030, nc18031, nc18032, 
        nc18033, nc18034, nc18035, nc18036, nc18037, nc18038, nc18039, 
        nc18040, nc18041, nc18042, nc18043, nc18044, nc18045, nc18046, 
        nc18047, nc18048, nc18049}), .DB_DETECT(\DB_DETECT[0][0] ), 
        .SB_CORRECT(\SB_CORRECT[0][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C9 (.A_DOUT({
        nc18050, nc18051, nc18052, nc18053, nc18054, nc18055, nc18056, 
        nc18057, nc18058, nc18059, nc18060, nc18061, nc18062, nc18063, 
        nc18064, nc18065, nc18066, nc18067, \R_DATA_TEMPR29[19] , 
        \R_DATA_TEMPR29[18] }), .B_DOUT({nc18068, nc18069, nc18070, 
        nc18071, nc18072, nc18073, nc18074, nc18075, nc18076, nc18077, 
        nc18078, nc18079, nc18080, nc18081, nc18082, nc18083, nc18084, 
        nc18085, nc18086, nc18087}), .DB_DETECT(\DB_DETECT[29][9] ), 
        .SB_CORRECT(\SB_CORRECT[29][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C11 (.A_DOUT({
        nc18088, nc18089, nc18090, nc18091, nc18092, nc18093, nc18094, 
        nc18095, nc18096, nc18097, nc18098, nc18099, nc18100, nc18101, 
        nc18102, nc18103, nc18104, nc18105, \R_DATA_TEMPR15[23] , 
        \R_DATA_TEMPR15[22] }), .B_DOUT({nc18106, nc18107, nc18108, 
        nc18109, nc18110, nc18111, nc18112, nc18113, nc18114, nc18115, 
        nc18116, nc18117, nc18118, nc18119, nc18120, nc18121, nc18122, 
        nc18123, nc18124, nc18125}), .DB_DETECT(\DB_DETECT[15][11] ), 
        .SB_CORRECT(\SB_CORRECT[15][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C7 (.A_DOUT({
        nc18126, nc18127, nc18128, nc18129, nc18130, nc18131, nc18132, 
        nc18133, nc18134, nc18135, nc18136, nc18137, nc18138, nc18139, 
        nc18140, nc18141, nc18142, nc18143, \R_DATA_TEMPR15[15] , 
        \R_DATA_TEMPR15[14] }), .B_DOUT({nc18144, nc18145, nc18146, 
        nc18147, nc18148, nc18149, nc18150, nc18151, nc18152, nc18153, 
        nc18154, nc18155, nc18156, nc18157, nc18158, nc18159, nc18160, 
        nc18161, nc18162, nc18163}), .DB_DETECT(\DB_DETECT[15][7] ), 
        .SB_CORRECT(\SB_CORRECT[15][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C2 (.A_DOUT({nc18164, 
        nc18165, nc18166, nc18167, nc18168, nc18169, nc18170, nc18171, 
        nc18172, nc18173, nc18174, nc18175, nc18176, nc18177, nc18178, 
        nc18179, nc18180, nc18181, \R_DATA_TEMPR6[5] , 
        \R_DATA_TEMPR6[4] }), .B_DOUT({nc18182, nc18183, nc18184, 
        nc18185, nc18186, nc18187, nc18188, nc18189, nc18190, nc18191, 
        nc18192, nc18193, nc18194, nc18195, nc18196, nc18197, nc18198, 
        nc18199, nc18200, nc18201}), .DB_DETECT(\DB_DETECT[6][2] ), 
        .SB_CORRECT(\SB_CORRECT[6][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_352 (.A(\R_DATA_TEMPR24[35] ), .B(\R_DATA_TEMPR25[35] ), 
        .C(\R_DATA_TEMPR26[35] ), .D(\R_DATA_TEMPR27[35] ), .Y(
        OR4_352_Y));
    OR4 OR4_15 (.A(OR4_183_Y), .B(OR2_18_Y), .C(\R_DATA_TEMPR22[38] ), 
        .D(\R_DATA_TEMPR23[38] ), .Y(OR4_15_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C2 (.A_DOUT({
        nc18202, nc18203, nc18204, nc18205, nc18206, nc18207, nc18208, 
        nc18209, nc18210, nc18211, nc18212, nc18213, nc18214, nc18215, 
        nc18216, nc18217, nc18218, nc18219, \R_DATA_TEMPR28[5] , 
        \R_DATA_TEMPR28[4] }), .B_DOUT({nc18220, nc18221, nc18222, 
        nc18223, nc18224, nc18225, nc18226, nc18227, nc18228, nc18229, 
        nc18230, nc18231, nc18232, nc18233, nc18234, nc18235, nc18236, 
        nc18237, nc18238, nc18239}), .DB_DETECT(\DB_DETECT[28][2] ), 
        .SB_CORRECT(\SB_CORRECT[28][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[28][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[3]  (.A(CFG2_0_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[3] ));
    OR4 OR4_281 (.A(\R_DATA_TEMPR16[37] ), .B(\R_DATA_TEMPR17[37] ), 
        .C(\R_DATA_TEMPR18[37] ), .D(\R_DATA_TEMPR19[37] ), .Y(
        OR4_281_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C10 (.A_DOUT({
        nc18240, nc18241, nc18242, nc18243, nc18244, nc18245, nc18246, 
        nc18247, nc18248, nc18249, nc18250, nc18251, nc18252, nc18253, 
        nc18254, nc18255, nc18256, nc18257, \R_DATA_TEMPR17[21] , 
        \R_DATA_TEMPR17[20] }), .B_DOUT({nc18258, nc18259, nc18260, 
        nc18261, nc18262, nc18263, nc18264, nc18265, nc18266, nc18267, 
        nc18268, nc18269, nc18270, nc18271, nc18272, nc18273, nc18274, 
        nc18275, nc18276, nc18277}), .DB_DETECT(\DB_DETECT[17][10] ), 
        .SB_CORRECT(\SB_CORRECT[17][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C3 (.A_DOUT({
        nc18278, nc18279, nc18280, nc18281, nc18282, nc18283, nc18284, 
        nc18285, nc18286, nc18287, nc18288, nc18289, nc18290, nc18291, 
        nc18292, nc18293, nc18294, nc18295, \R_DATA_TEMPR16[7] , 
        \R_DATA_TEMPR16[6] }), .B_DOUT({nc18296, nc18297, nc18298, 
        nc18299, nc18300, nc18301, nc18302, nc18303, nc18304, nc18305, 
        nc18306, nc18307, nc18308, nc18309, nc18310, nc18311, nc18312, 
        nc18313, nc18314, nc18315}), .DB_DETECT(\DB_DETECT[16][3] ), 
        .SB_CORRECT(\SB_CORRECT[16][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_326 (.A(\R_DATA_TEMPR0[1] ), .B(\R_DATA_TEMPR1[1] ), .C(
        \R_DATA_TEMPR2[1] ), .D(\R_DATA_TEMPR3[1] ), .Y(OR4_326_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C14 (.A_DOUT({
        nc18316, nc18317, nc18318, nc18319, nc18320, nc18321, nc18322, 
        nc18323, nc18324, nc18325, nc18326, nc18327, nc18328, nc18329, 
        nc18330, nc18331, nc18332, nc18333, \R_DATA_TEMPR13[29] , 
        \R_DATA_TEMPR13[28] }), .B_DOUT({nc18334, nc18335, nc18336, 
        nc18337, nc18338, nc18339, nc18340, nc18341, nc18342, nc18343, 
        nc18344, nc18345, nc18346, nc18347, nc18348, nc18349, nc18350, 
        nc18351, nc18352, nc18353}), .DB_DETECT(\DB_DETECT[13][14] ), 
        .SB_CORRECT(\SB_CORRECT[13][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_194 (.A(\R_DATA_TEMPR12[38] ), .B(\R_DATA_TEMPR13[38] ), 
        .C(\R_DATA_TEMPR14[38] ), .D(\R_DATA_TEMPR15[38] ), .Y(
        OR4_194_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C15 (.A_DOUT({
        nc18354, nc18355, nc18356, nc18357, nc18358, nc18359, nc18360, 
        nc18361, nc18362, nc18363, nc18364, nc18365, nc18366, nc18367, 
        nc18368, nc18369, nc18370, nc18371, \R_DATA_TEMPR30[31] , 
        \R_DATA_TEMPR30[30] }), .B_DOUT({nc18372, nc18373, nc18374, 
        nc18375, nc18376, nc18377, nc18378, nc18379, nc18380, nc18381, 
        nc18382, nc18383, nc18384, nc18385, nc18386, nc18387, nc18388, 
        nc18389, nc18390, nc18391}), .DB_DETECT(\DB_DETECT[30][15] ), 
        .SB_CORRECT(\SB_CORRECT[30][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C15 (.A_DOUT({
        nc18392, nc18393, nc18394, nc18395, nc18396, nc18397, nc18398, 
        nc18399, nc18400, nc18401, nc18402, nc18403, nc18404, nc18405, 
        nc18406, nc18407, nc18408, nc18409, \R_DATA_TEMPR17[31] , 
        \R_DATA_TEMPR17[30] }), .B_DOUT({nc18410, nc18411, nc18412, 
        nc18413, nc18414, nc18415, nc18416, nc18417, nc18418, nc18419, 
        nc18420, nc18421, nc18422, nc18423, nc18424, nc18425, nc18426, 
        nc18427, nc18428, nc18429}), .DB_DETECT(\DB_DETECT[17][15] ), 
        .SB_CORRECT(\SB_CORRECT[17][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_93 (.A(\R_DATA_TEMPR12[23] ), .B(\R_DATA_TEMPR13[23] ), .C(
        \R_DATA_TEMPR14[23] ), .D(\R_DATA_TEMPR15[23] ), .Y(OR4_93_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C10 (.A_DOUT({
        nc18430, nc18431, nc18432, nc18433, nc18434, nc18435, nc18436, 
        nc18437, nc18438, nc18439, nc18440, nc18441, nc18442, nc18443, 
        nc18444, nc18445, nc18446, nc18447, \R_DATA_TEMPR8[21] , 
        \R_DATA_TEMPR8[20] }), .B_DOUT({nc18448, nc18449, nc18450, 
        nc18451, nc18452, nc18453, nc18454, nc18455, nc18456, nc18457, 
        nc18458, nc18459, nc18460, nc18461, nc18462, nc18463, nc18464, 
        nc18465, nc18466, nc18467}), .DB_DETECT(\DB_DETECT[8][10] ), 
        .SB_CORRECT(\SB_CORRECT[8][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_309 (.A(\R_DATA_TEMPR16[14] ), .B(\R_DATA_TEMPR17[14] ), 
        .C(\R_DATA_TEMPR18[14] ), .D(\R_DATA_TEMPR19[14] ), .Y(
        OR4_309_Y));
    OR4 OR4_24 (.A(\R_DATA_TEMPR8[1] ), .B(\R_DATA_TEMPR9[1] ), .C(
        \R_DATA_TEMPR10[1] ), .D(\R_DATA_TEMPR11[1] ), .Y(OR4_24_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C3 (.A_DOUT({
        nc18468, nc18469, nc18470, nc18471, nc18472, nc18473, nc18474, 
        nc18475, nc18476, nc18477, nc18478, nc18479, nc18480, nc18481, 
        nc18482, nc18483, nc18484, nc18485, \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR10[6] }), .B_DOUT({nc18486, nc18487, nc18488, 
        nc18489, nc18490, nc18491, nc18492, nc18493, nc18494, nc18495, 
        nc18496, nc18497, nc18498, nc18499, nc18500, nc18501, nc18502, 
        nc18503, nc18504, nc18505}), .DB_DETECT(\DB_DETECT[10][3] ), 
        .SB_CORRECT(\SB_CORRECT[10][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C3 (.A_DOUT({
        nc18506, nc18507, nc18508, nc18509, nc18510, nc18511, nc18512, 
        nc18513, nc18514, nc18515, nc18516, nc18517, nc18518, nc18519, 
        nc18520, nc18521, nc18522, nc18523, \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR13[6] }), .B_DOUT({nc18524, nc18525, nc18526, 
        nc18527, nc18528, nc18529, nc18530, nc18531, nc18532, nc18533, 
        nc18534, nc18535, nc18536, nc18537, nc18538, nc18539, nc18540, 
        nc18541, nc18542, nc18543}), .DB_DETECT(\DB_DETECT[13][3] ), 
        .SB_CORRECT(\SB_CORRECT[13][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_8 (.A(\R_DATA_TEMPR8[24] ), .B(\R_DATA_TEMPR9[24] ), .C(
        \R_DATA_TEMPR10[24] ), .D(\R_DATA_TEMPR11[24] ), .Y(OR4_8_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C19 (.A_DOUT({
        nc18544, nc18545, nc18546, nc18547, nc18548, nc18549, nc18550, 
        nc18551, nc18552, nc18553, nc18554, nc18555, nc18556, nc18557, 
        nc18558, nc18559, nc18560, nc18561, \R_DATA_TEMPR18[39] , 
        \R_DATA_TEMPR18[38] }), .B_DOUT({nc18562, nc18563, nc18564, 
        nc18565, nc18566, nc18567, nc18568, nc18569, nc18570, nc18571, 
        nc18572, nc18573, nc18574, nc18575, nc18576, nc18577, nc18578, 
        nc18579, nc18580, nc18581}), .DB_DETECT(\DB_DETECT[18][19] ), 
        .SB_CORRECT(\SB_CORRECT[18][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_250 (.A(\R_DATA_TEMPR12[17] ), .B(\R_DATA_TEMPR13[17] ), 
        .C(\R_DATA_TEMPR14[17] ), .D(\R_DATA_TEMPR15[17] ), .Y(
        OR4_250_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C18 (.A_DOUT({
        nc18582, nc18583, nc18584, nc18585, nc18586, nc18587, nc18588, 
        nc18589, nc18590, nc18591, nc18592, nc18593, nc18594, nc18595, 
        nc18596, nc18597, nc18598, nc18599, \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR4[36] }), .B_DOUT({nc18600, nc18601, nc18602, 
        nc18603, nc18604, nc18605, nc18606, nc18607, nc18608, nc18609, 
        nc18610, nc18611, nc18612, nc18613, nc18614, nc18615, nc18616, 
        nc18617, nc18618, nc18619}), .DB_DETECT(\DB_DETECT[4][18] ), 
        .SB_CORRECT(\SB_CORRECT[4][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C9 (.A_DOUT({
        nc18620, nc18621, nc18622, nc18623, nc18624, nc18625, nc18626, 
        nc18627, nc18628, nc18629, nc18630, nc18631, nc18632, nc18633, 
        nc18634, nc18635, nc18636, nc18637, \R_DATA_TEMPR28[19] , 
        \R_DATA_TEMPR28[18] }), .B_DOUT({nc18638, nc18639, nc18640, 
        nc18641, nc18642, nc18643, nc18644, nc18645, nc18646, nc18647, 
        nc18648, nc18649, nc18650, nc18651, nc18652, nc18653, nc18654, 
        nc18655, nc18656, nc18657}), .DB_DETECT(\DB_DETECT[28][9] ), 
        .SB_CORRECT(\SB_CORRECT[28][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[28][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_334 (.A(OR4_209_Y), .B(OR2_34_Y), .C(\R_DATA_TEMPR22[1] ), 
        .D(\R_DATA_TEMPR23[1] ), .Y(OR4_334_Y));
    OR2 OR2_4 (.A(\R_DATA_TEMPR20[10] ), .B(\R_DATA_TEMPR21[10] ), .Y(
        OR2_4_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C2 (.A_DOUT({nc18658, 
        nc18659, nc18660, nc18661, nc18662, nc18663, nc18664, nc18665, 
        nc18666, nc18667, nc18668, nc18669, nc18670, nc18671, nc18672, 
        nc18673, nc18674, nc18675, \R_DATA_TEMPR9[5] , 
        \R_DATA_TEMPR9[4] }), .B_DOUT({nc18676, nc18677, nc18678, 
        nc18679, nc18680, nc18681, nc18682, nc18683, nc18684, nc18685, 
        nc18686, nc18687, nc18688, nc18689, nc18690, nc18691, nc18692, 
        nc18693, nc18694, nc18695}), .DB_DETECT(\DB_DETECT[9][2] ), 
        .SB_CORRECT(\SB_CORRECT[9][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C16 (.A_DOUT({
        nc18696, nc18697, nc18698, nc18699, nc18700, nc18701, nc18702, 
        nc18703, nc18704, nc18705, nc18706, nc18707, nc18708, nc18709, 
        nc18710, nc18711, nc18712, nc18713, \R_DATA_TEMPR0[33] , 
        \R_DATA_TEMPR0[32] }), .B_DOUT({nc18714, nc18715, nc18716, 
        nc18717, nc18718, nc18719, nc18720, nc18721, nc18722, nc18723, 
        nc18724, nc18725, nc18726, nc18727, nc18728, nc18729, nc18730, 
        nc18731, nc18732, nc18733}), .DB_DETECT(\DB_DETECT[0][16] ), 
        .SB_CORRECT(\SB_CORRECT[0][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C2 (.A_DOUT({
        nc18734, nc18735, nc18736, nc18737, nc18738, nc18739, nc18740, 
        nc18741, nc18742, nc18743, nc18744, nc18745, nc18746, nc18747, 
        nc18748, nc18749, nc18750, nc18751, \R_DATA_TEMPR11[5] , 
        \R_DATA_TEMPR11[4] }), .B_DOUT({nc18752, nc18753, nc18754, 
        nc18755, nc18756, nc18757, nc18758, nc18759, nc18760, nc18761, 
        nc18762, nc18763, nc18764, nc18765, nc18766, nc18767, nc18768, 
        nc18769, nc18770, nc18771}), .DB_DETECT(\DB_DETECT[11][2] ), 
        .SB_CORRECT(\SB_CORRECT[11][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_131 (.A(\R_DATA_TEMPR4[28] ), .B(\R_DATA_TEMPR5[28] ), .C(
        \R_DATA_TEMPR6[28] ), .D(\R_DATA_TEMPR7[28] ), .Y(OR4_131_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C3 (.A_DOUT({nc18772, 
        nc18773, nc18774, nc18775, nc18776, nc18777, nc18778, nc18779, 
        nc18780, nc18781, nc18782, nc18783, nc18784, nc18785, nc18786, 
        nc18787, nc18788, nc18789, \R_DATA_TEMPR1[7] , 
        \R_DATA_TEMPR1[6] }), .B_DOUT({nc18790, nc18791, nc18792, 
        nc18793, nc18794, nc18795, nc18796, nc18797, nc18798, nc18799, 
        nc18800, nc18801, nc18802, nc18803, nc18804, nc18805, nc18806, 
        nc18807, nc18808, nc18809}), .DB_DETECT(\DB_DETECT[1][3] ), 
        .SB_CORRECT(\SB_CORRECT[1][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C18 (.A_DOUT({
        nc18810, nc18811, nc18812, nc18813, nc18814, nc18815, nc18816, 
        nc18817, nc18818, nc18819, nc18820, nc18821, nc18822, nc18823, 
        nc18824, nc18825, nc18826, nc18827, \R_DATA_TEMPR19[37] , 
        \R_DATA_TEMPR19[36] }), .B_DOUT({nc18828, nc18829, nc18830, 
        nc18831, nc18832, nc18833, nc18834, nc18835, nc18836, nc18837, 
        nc18838, nc18839, nc18840, nc18841, nc18842, nc18843, nc18844, 
        nc18845, nc18846, nc18847}), .DB_DETECT(\DB_DETECT[19][18] ), 
        .SB_CORRECT(\SB_CORRECT[19][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C19 (.A_DOUT({
        nc18848, nc18849, nc18850, nc18851, nc18852, nc18853, nc18854, 
        nc18855, nc18856, nc18857, nc18858, nc18859, nc18860, nc18861, 
        nc18862, nc18863, nc18864, nc18865, \R_DATA_TEMPR9[39] , 
        \R_DATA_TEMPR9[38] }), .B_DOUT({nc18866, nc18867, nc18868, 
        nc18869, nc18870, nc18871, nc18872, nc18873, nc18874, nc18875, 
        nc18876, nc18877, nc18878, nc18879, nc18880, nc18881, nc18882, 
        nc18883, nc18884, nc18885}), .DB_DETECT(\DB_DETECT[9][19] ), 
        .SB_CORRECT(\SB_CORRECT[9][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[39]  (.A(OR4_193_Y), .B(OR4_122_Y), .C(OR4_95_Y), 
        .D(OR4_22_Y), .Y(R_DATA[39]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C9 (.A_DOUT({
        nc18886, nc18887, nc18888, nc18889, nc18890, nc18891, nc18892, 
        nc18893, nc18894, nc18895, nc18896, nc18897, nc18898, nc18899, 
        nc18900, nc18901, nc18902, nc18903, \R_DATA_TEMPR22[19] , 
        \R_DATA_TEMPR22[18] }), .B_DOUT({nc18904, nc18905, nc18906, 
        nc18907, nc18908, nc18909, nc18910, nc18911, nc18912, nc18913, 
        nc18914, nc18915, nc18916, nc18917, nc18918, nc18919, nc18920, 
        nc18921, nc18922, nc18923}), .DB_DETECT(\DB_DETECT[22][9] ), 
        .SB_CORRECT(\SB_CORRECT[22][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_256 (.A(OR4_324_Y), .B(OR4_169_Y), .C(OR4_247_Y), .D(
        OR4_72_Y), .Y(OR4_256_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C9 (.A_DOUT({
        nc18924, nc18925, nc18926, nc18927, nc18928, nc18929, nc18930, 
        nc18931, nc18932, nc18933, nc18934, nc18935, nc18936, nc18937, 
        nc18938, nc18939, nc18940, nc18941, \R_DATA_TEMPR15[19] , 
        \R_DATA_TEMPR15[18] }), .B_DOUT({nc18942, nc18943, nc18944, 
        nc18945, nc18946, nc18947, nc18948, nc18949, nc18950, nc18951, 
        nc18952, nc18953, nc18954, nc18955, nc18956, nc18957, nc18958, 
        nc18959, nc18960, nc18961}), .DB_DETECT(\DB_DETECT[15][9] ), 
        .SB_CORRECT(\SB_CORRECT[15][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_0 (.A(\R_DATA_TEMPR20[12] ), .B(\R_DATA_TEMPR21[12] ), .Y(
        OR2_0_Y));
    OR4 OR4_75 (.A(\R_DATA_TEMPR4[8] ), .B(\R_DATA_TEMPR5[8] ), .C(
        \R_DATA_TEMPR6[8] ), .D(\R_DATA_TEMPR7[8] ), .Y(OR4_75_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C9 (.A_DOUT({nc18962, 
        nc18963, nc18964, nc18965, nc18966, nc18967, nc18968, nc18969, 
        nc18970, nc18971, nc18972, nc18973, nc18974, nc18975, nc18976, 
        nc18977, nc18978, nc18979, \R_DATA_TEMPR4[19] , 
        \R_DATA_TEMPR4[18] }), .B_DOUT({nc18980, nc18981, nc18982, 
        nc18983, nc18984, nc18985, nc18986, nc18987, nc18988, nc18989, 
        nc18990, nc18991, nc18992, nc18993, nc18994, nc18995, nc18996, 
        nc18997, nc18998, nc18999}), .DB_DETECT(\DB_DETECT[4][9] ), 
        .SB_CORRECT(\SB_CORRECT[4][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_6 (.A(\R_DATA_TEMPR20[32] ), .B(\R_DATA_TEMPR21[32] ), .Y(
        OR2_6_Y));
    OR4 OR4_91 (.A(\R_DATA_TEMPR16[16] ), .B(\R_DATA_TEMPR17[16] ), .C(
        \R_DATA_TEMPR18[16] ), .D(\R_DATA_TEMPR19[16] ), .Y(OR4_91_Y));
    OR4 OR4_124 (.A(\R_DATA_TEMPR28[32] ), .B(\R_DATA_TEMPR29[32] ), 
        .C(\R_DATA_TEMPR30[32] ), .D(\R_DATA_TEMPR31[32] ), .Y(
        OR4_124_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0 (.A_DOUT({nc19000, 
        nc19001, nc19002, nc19003, nc19004, nc19005, nc19006, nc19007, 
        nc19008, nc19009, nc19010, nc19011, nc19012, nc19013, nc19014, 
        nc19015, nc19016, nc19017, \R_DATA_TEMPR6[1] , 
        \R_DATA_TEMPR6[0] }), .B_DOUT({nc19018, nc19019, nc19020, 
        nc19021, nc19022, nc19023, nc19024, nc19025, nc19026, nc19027, 
        nc19028, nc19029, nc19030, nc19031, nc19032, nc19033, nc19034, 
        nc19035, nc19036, nc19037}), .DB_DETECT(\DB_DETECT[6][0] ), 
        .SB_CORRECT(\SB_CORRECT[6][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C9 (.A_DOUT({
        nc19038, nc19039, nc19040, nc19041, nc19042, nc19043, nc19044, 
        nc19045, nc19046, nc19047, nc19048, nc19049, nc19050, nc19051, 
        nc19052, nc19053, nc19054, nc19055, \R_DATA_TEMPR11[19] , 
        \R_DATA_TEMPR11[18] }), .B_DOUT({nc19056, nc19057, nc19058, 
        nc19059, nc19060, nc19061, nc19062, nc19063, nc19064, nc19065, 
        nc19066, nc19067, nc19068, nc19069, nc19070, nc19071, nc19072, 
        nc19073, nc19074, nc19075}), .DB_DETECT(\DB_DETECT[11][9] ), 
        .SB_CORRECT(\SB_CORRECT[11][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_3 (.A(\R_DATA_TEMPR20[9] ), .B(\R_DATA_TEMPR21[9] ), .Y(
        OR2_3_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[5]  (.A(CFG2_2_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[5] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C10 (.A_DOUT({
        nc19076, nc19077, nc19078, nc19079, nc19080, nc19081, nc19082, 
        nc19083, nc19084, nc19085, nc19086, nc19087, nc19088, nc19089, 
        nc19090, nc19091, nc19092, nc19093, \R_DATA_TEMPR12[21] , 
        \R_DATA_TEMPR12[20] }), .B_DOUT({nc19094, nc19095, nc19096, 
        nc19097, nc19098, nc19099, nc19100, nc19101, nc19102, nc19103, 
        nc19104, nc19105, nc19106, nc19107, nc19108, nc19109, nc19110, 
        nc19111, nc19112, nc19113}), .DB_DETECT(\DB_DETECT[12][10] ), 
        .SB_CORRECT(\SB_CORRECT[12][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C4 (.A_DOUT({nc19114, 
        nc19115, nc19116, nc19117, nc19118, nc19119, nc19120, nc19121, 
        nc19122, nc19123, nc19124, nc19125, nc19126, nc19127, nc19128, 
        nc19129, nc19130, nc19131, \R_DATA_TEMPR0[9] , 
        \R_DATA_TEMPR0[8] }), .B_DOUT({nc19132, nc19133, nc19134, 
        nc19135, nc19136, nc19137, nc19138, nc19139, nc19140, nc19141, 
        nc19142, nc19143, nc19144, nc19145, nc19146, nc19147, nc19148, 
        nc19149, nc19150, nc19151}), .DB_DETECT(\DB_DETECT[0][4] ), 
        .SB_CORRECT(\SB_CORRECT[0][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C14 (.A_DOUT({
        nc19152, nc19153, nc19154, nc19155, nc19156, nc19157, nc19158, 
        nc19159, nc19160, nc19161, nc19162, nc19163, nc19164, nc19165, 
        nc19166, nc19167, nc19168, nc19169, \R_DATA_TEMPR3[29] , 
        \R_DATA_TEMPR3[28] }), .B_DOUT({nc19170, nc19171, nc19172, 
        nc19173, nc19174, nc19175, nc19176, nc19177, nc19178, nc19179, 
        nc19180, nc19181, nc19182, nc19183, nc19184, nc19185, nc19186, 
        nc19187, nc19188, nc19189}), .DB_DETECT(\DB_DETECT[3][14] ), 
        .SB_CORRECT(\SB_CORRECT[3][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C15 (.A_DOUT({
        nc19190, nc19191, nc19192, nc19193, nc19194, nc19195, nc19196, 
        nc19197, nc19198, nc19199, nc19200, nc19201, nc19202, nc19203, 
        nc19204, nc19205, nc19206, nc19207, \R_DATA_TEMPR12[31] , 
        \R_DATA_TEMPR12[30] }), .B_DOUT({nc19208, nc19209, nc19210, 
        nc19211, nc19212, nc19213, nc19214, nc19215, nc19216, nc19217, 
        nc19218, nc19219, nc19220, nc19221, nc19222, nc19223, nc19224, 
        nc19225, nc19226, nc19227}), .DB_DETECT(\DB_DETECT[12][15] ), 
        .SB_CORRECT(\SB_CORRECT[12][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C8 (.A_DOUT({
        nc19228, nc19229, nc19230, nc19231, nc19232, nc19233, nc19234, 
        nc19235, nc19236, nc19237, nc19238, nc19239, nc19240, nc19241, 
        nc19242, nc19243, nc19244, nc19245, \R_DATA_TEMPR24[17] , 
        \R_DATA_TEMPR24[16] }), .B_DOUT({nc19246, nc19247, nc19248, 
        nc19249, nc19250, nc19251, nc19252, nc19253, nc19254, nc19255, 
        nc19256, nc19257, nc19258, nc19259, nc19260, nc19261, nc19262, 
        nc19263, nc19264, nc19265}), .DB_DETECT(\DB_DETECT[24][8] ), 
        .SB_CORRECT(\SB_CORRECT[24][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[7]  (.A(CFG2_0_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[7] ));
    OR4 OR4_314 (.A(\R_DATA_TEMPR0[38] ), .B(\R_DATA_TEMPR1[38] ), .C(
        \R_DATA_TEMPR2[38] ), .D(\R_DATA_TEMPR3[38] ), .Y(OR4_314_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C4 (.A_DOUT({
        nc19266, nc19267, nc19268, nc19269, nc19270, nc19271, nc19272, 
        nc19273, nc19274, nc19275, nc19276, nc19277, nc19278, nc19279, 
        nc19280, nc19281, nc19282, nc19283, \R_DATA_TEMPR27[9] , 
        \R_DATA_TEMPR27[8] }), .B_DOUT({nc19284, nc19285, nc19286, 
        nc19287, nc19288, nc19289, nc19290, nc19291, nc19292, nc19293, 
        nc19294, nc19295, nc19296, nc19297, nc19298, nc19299, nc19300, 
        nc19301, nc19302, nc19303}), .DB_DETECT(\DB_DETECT[27][4] ), 
        .SB_CORRECT(\SB_CORRECT[27][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0 (.A_DOUT({
        nc19304, nc19305, nc19306, nc19307, nc19308, nc19309, nc19310, 
        nc19311, nc19312, nc19313, nc19314, nc19315, nc19316, nc19317, 
        nc19318, nc19319, nc19320, nc19321, \R_DATA_TEMPR28[1] , 
        \R_DATA_TEMPR28[0] }), .B_DOUT({nc19322, nc19323, nc19324, 
        nc19325, nc19326, nc19327, nc19328, nc19329, nc19330, nc19331, 
        nc19332, nc19333, nc19334, nc19335, nc19336, nc19337, nc19338, 
        nc19339, nc19340, nc19341}), .DB_DETECT(\DB_DETECT[28][0] ), 
        .SB_CORRECT(\SB_CORRECT[28][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[28][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C1 (.A_DOUT({
        nc19342, nc19343, nc19344, nc19345, nc19346, nc19347, nc19348, 
        nc19349, nc19350, nc19351, nc19352, nc19353, nc19354, nc19355, 
        nc19356, nc19357, nc19358, nc19359, \R_DATA_TEMPR28[3] , 
        \R_DATA_TEMPR28[2] }), .B_DOUT({nc19360, nc19361, nc19362, 
        nc19363, nc19364, nc19365, nc19366, nc19367, nc19368, nc19369, 
        nc19370, nc19371, nc19372, nc19373, nc19374, nc19375, nc19376, 
        nc19377, nc19378, nc19379}), .DB_DETECT(\DB_DETECT[28][1] ), 
        .SB_CORRECT(\SB_CORRECT[28][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[28][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C3 (.A_DOUT({
        nc19380, nc19381, nc19382, nc19383, nc19384, nc19385, nc19386, 
        nc19387, nc19388, nc19389, nc19390, nc19391, nc19392, nc19393, 
        nc19394, nc19395, nc19396, nc19397, \R_DATA_TEMPR19[7] , 
        \R_DATA_TEMPR19[6] }), .B_DOUT({nc19398, nc19399, nc19400, 
        nc19401, nc19402, nc19403, nc19404, nc19405, nc19406, nc19407, 
        nc19408, nc19409, nc19410, nc19411, nc19412, nc19413, nc19414, 
        nc19415, nc19416, nc19417}), .DB_DETECT(\DB_DETECT[19][3] ), 
        .SB_CORRECT(\SB_CORRECT[19][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C2 (.A_DOUT({
        nc19418, nc19419, nc19420, nc19421, nc19422, nc19423, nc19424, 
        nc19425, nc19426, nc19427, nc19428, nc19429, nc19430, nc19431, 
        nc19432, nc19433, nc19434, nc19435, \R_DATA_TEMPR30[5] , 
        \R_DATA_TEMPR30[4] }), .B_DOUT({nc19436, nc19437, nc19438, 
        nc19439, nc19440, nc19441, nc19442, nc19443, nc19444, nc19445, 
        nc19446, nc19447, nc19448, nc19449, nc19450, nc19451, nc19452, 
        nc19453, nc19454, nc19455}), .DB_DETECT(\DB_DETECT[30][2] ), 
        .SB_CORRECT(\SB_CORRECT[30][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[30][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_43 (.A(\R_DATA_TEMPR0[6] ), .B(\R_DATA_TEMPR1[6] ), .C(
        \R_DATA_TEMPR2[6] ), .D(\R_DATA_TEMPR3[6] ), .Y(OR4_43_Y));
    INV \INVBLKX0[0]  (.A(W_ADDR[13]), .Y(\BLKX0[0] ));
    OR2 OR2_26 (.A(\R_DATA_TEMPR20[24] ), .B(\R_DATA_TEMPR21[24] ), .Y(
        OR2_26_Y));
    OR4 OR4_111 (.A(\R_DATA_TEMPR4[4] ), .B(\R_DATA_TEMPR5[4] ), .C(
        \R_DATA_TEMPR6[4] ), .D(\R_DATA_TEMPR7[4] ), .Y(OR4_111_Y));
    OR4 OR4_59 (.A(\R_DATA_TEMPR0[25] ), .B(\R_DATA_TEMPR1[25] ), .C(
        \R_DATA_TEMPR2[25] ), .D(\R_DATA_TEMPR3[25] ), .Y(OR4_59_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0 (.A_DOUT({
        nc19456, nc19457, nc19458, nc19459, nc19460, nc19461, nc19462, 
        nc19463, nc19464, nc19465, nc19466, nc19467, nc19468, nc19469, 
        nc19470, nc19471, nc19472, nc19473, \R_DATA_TEMPR14[1] , 
        \R_DATA_TEMPR14[0] }), .B_DOUT({nc19474, nc19475, nc19476, 
        nc19477, nc19478, nc19479, nc19480, nc19481, nc19482, nc19483, 
        nc19484, nc19485, nc19486, nc19487, nc19488, nc19489, nc19490, 
        nc19491, nc19492, nc19493}), .DB_DETECT(\DB_DETECT[14][0] ), 
        .SB_CORRECT(\SB_CORRECT[14][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C14 (.A_DOUT({
        nc19494, nc19495, nc19496, nc19497, nc19498, nc19499, nc19500, 
        nc19501, nc19502, nc19503, nc19504, nc19505, nc19506, nc19507, 
        nc19508, nc19509, nc19510, nc19511, \R_DATA_TEMPR10[29] , 
        \R_DATA_TEMPR10[28] }), .B_DOUT({nc19512, nc19513, nc19514, 
        nc19515, nc19516, nc19517, nc19518, nc19519, nc19520, nc19521, 
        nc19522, nc19523, nc19524, nc19525, nc19526, nc19527, nc19528, 
        nc19529, nc19530, nc19531}), .DB_DETECT(\DB_DETECT[10][14] ), 
        .SB_CORRECT(\SB_CORRECT[10][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C1 (.A_DOUT({
        nc19532, nc19533, nc19534, nc19535, nc19536, nc19537, nc19538, 
        nc19539, nc19540, nc19541, nc19542, nc19543, nc19544, nc19545, 
        nc19546, nc19547, nc19548, nc19549, \R_DATA_TEMPR19[3] , 
        \R_DATA_TEMPR19[2] }), .B_DOUT({nc19550, nc19551, nc19552, 
        nc19553, nc19554, nc19555, nc19556, nc19557, nc19558, nc19559, 
        nc19560, nc19561, nc19562, nc19563, nc19564, nc19565, nc19566, 
        nc19567, nc19568, nc19569}), .DB_DETECT(\DB_DETECT[19][1] ), 
        .SB_CORRECT(\SB_CORRECT[19][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C19 (.A_DOUT({
        nc19570, nc19571, nc19572, nc19573, nc19574, nc19575, nc19576, 
        nc19577, nc19578, nc19579, nc19580, nc19581, nc19582, nc19583, 
        nc19584, nc19585, nc19586, nc19587, \R_DATA_TEMPR23[39] , 
        \R_DATA_TEMPR23[38] }), .B_DOUT({nc19588, nc19589, nc19590, 
        nc19591, nc19592, nc19593, nc19594, nc19595, nc19596, nc19597, 
        nc19598, nc19599, nc19600, nc19601, nc19602, nc19603, nc19604, 
        nc19605, nc19606, nc19607}), .DB_DETECT(\DB_DETECT[23][19] ), 
        .SB_CORRECT(\SB_CORRECT[23][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_263 (.A(\R_DATA_TEMPR24[15] ), .B(\R_DATA_TEMPR25[15] ), 
        .C(\R_DATA_TEMPR26[15] ), .D(\R_DATA_TEMPR27[15] ), .Y(
        OR4_263_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C9 (.A_DOUT({
        nc19608, nc19609, nc19610, nc19611, nc19612, nc19613, nc19614, 
        nc19615, nc19616, nc19617, nc19618, nc19619, nc19620, nc19621, 
        nc19622, nc19623, nc19624, nc19625, \R_DATA_TEMPR23[19] , 
        \R_DATA_TEMPR23[18] }), .B_DOUT({nc19626, nc19627, nc19628, 
        nc19629, nc19630, nc19631, nc19632, nc19633, nc19634, nc19635, 
        nc19636, nc19637, nc19638, nc19639, nc19640, nc19641, nc19642, 
        nc19643, nc19644, nc19645}), .DB_DETECT(\DB_DETECT[23][9] ), 
        .SB_CORRECT(\SB_CORRECT[23][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C3 (.A_DOUT({nc19646, 
        nc19647, nc19648, nc19649, nc19650, nc19651, nc19652, nc19653, 
        nc19654, nc19655, nc19656, nc19657, nc19658, nc19659, nc19660, 
        nc19661, nc19662, nc19663, \R_DATA_TEMPR4[7] , 
        \R_DATA_TEMPR4[6] }), .B_DOUT({nc19664, nc19665, nc19666, 
        nc19667, nc19668, nc19669, nc19670, nc19671, nc19672, nc19673, 
        nc19674, nc19675, nc19676, nc19677, nc19678, nc19679, nc19680, 
        nc19681, nc19682, nc19683}), .DB_DETECT(\DB_DETECT[4][3] ), 
        .SB_CORRECT(\SB_CORRECT[4][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C2 (.A_DOUT({nc19684, 
        nc19685, nc19686, nc19687, nc19688, nc19689, nc19690, nc19691, 
        nc19692, nc19693, nc19694, nc19695, nc19696, nc19697, nc19698, 
        nc19699, nc19700, nc19701, \R_DATA_TEMPR5[5] , 
        \R_DATA_TEMPR5[4] }), .B_DOUT({nc19702, nc19703, nc19704, 
        nc19705, nc19706, nc19707, nc19708, nc19709, nc19710, nc19711, 
        nc19712, nc19713, nc19714, nc19715, nc19716, nc19717, nc19718, 
        nc19719, nc19720, nc19721}), .DB_DETECT(\DB_DETECT[5][2] ), 
        .SB_CORRECT(\SB_CORRECT[5][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C5 (.A_DOUT({nc19722, 
        nc19723, nc19724, nc19725, nc19726, nc19727, nc19728, nc19729, 
        nc19730, nc19731, nc19732, nc19733, nc19734, nc19735, nc19736, 
        nc19737, nc19738, nc19739, \R_DATA_TEMPR4[11] , 
        \R_DATA_TEMPR4[10] }), .B_DOUT({nc19740, nc19741, nc19742, 
        nc19743, nc19744, nc19745, nc19746, nc19747, nc19748, nc19749, 
        nc19750, nc19751, nc19752, nc19753, nc19754, nc19755, nc19756, 
        nc19757, nc19758, nc19759}), .DB_DETECT(\DB_DETECT[4][5] ), 
        .SB_CORRECT(\SB_CORRECT[4][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C8 (.A_DOUT({
        nc19760, nc19761, nc19762, nc19763, nc19764, nc19765, nc19766, 
        nc19767, nc19768, nc19769, nc19770, nc19771, nc19772, nc19773, 
        nc19774, nc19775, nc19776, nc19777, \R_DATA_TEMPR11[17] , 
        \R_DATA_TEMPR11[16] }), .B_DOUT({nc19778, nc19779, nc19780, 
        nc19781, nc19782, nc19783, nc19784, nc19785, nc19786, nc19787, 
        nc19788, nc19789, nc19790, nc19791, nc19792, nc19793, nc19794, 
        nc19795, nc19796, nc19797}), .DB_DETECT(\DB_DETECT[11][8] ), 
        .SB_CORRECT(\SB_CORRECT[11][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[0]  (.A(OR4_297_Y), .B(OR4_337_Y), .C(OR4_220_Y), 
        .D(OR4_293_Y), .Y(R_DATA[0]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C6 (.A_DOUT({nc19798, 
        nc19799, nc19800, nc19801, nc19802, nc19803, nc19804, nc19805, 
        nc19806, nc19807, nc19808, nc19809, nc19810, nc19811, nc19812, 
        nc19813, nc19814, nc19815, \R_DATA_TEMPR9[13] , 
        \R_DATA_TEMPR9[12] }), .B_DOUT({nc19816, nc19817, nc19818, 
        nc19819, nc19820, nc19821, nc19822, nc19823, nc19824, nc19825, 
        nc19826, nc19827, nc19828, nc19829, nc19830, nc19831, nc19832, 
        nc19833, nc19834, nc19835}), .DB_DETECT(\DB_DETECT[9][6] ), 
        .SB_CORRECT(\SB_CORRECT[9][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C2 (.A_DOUT({
        nc19836, nc19837, nc19838, nc19839, nc19840, nc19841, nc19842, 
        nc19843, nc19844, nc19845, nc19846, nc19847, nc19848, nc19849, 
        nc19850, nc19851, nc19852, nc19853, \R_DATA_TEMPR24[5] , 
        \R_DATA_TEMPR24[4] }), .B_DOUT({nc19854, nc19855, nc19856, 
        nc19857, nc19858, nc19859, nc19860, nc19861, nc19862, nc19863, 
        nc19864, nc19865, nc19866, nc19867, nc19868, nc19869, nc19870, 
        nc19871, nc19872, nc19873}), .DB_DETECT(\DB_DETECT[24][2] ), 
        .SB_CORRECT(\SB_CORRECT[24][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_19 (.A(\R_DATA_TEMPR4[37] ), .B(\R_DATA_TEMPR5[37] ), .C(
        \R_DATA_TEMPR6[37] ), .D(\R_DATA_TEMPR7[37] ), .Y(OR4_19_Y));
    OR4 OR4_333 (.A(\R_DATA_TEMPR8[36] ), .B(\R_DATA_TEMPR9[36] ), .C(
        \R_DATA_TEMPR10[36] ), .D(\R_DATA_TEMPR11[36] ), .Y(OR4_333_Y));
    OR4 OR4_41 (.A(OR4_116_Y), .B(OR4_315_Y), .C(OR4_197_Y), .D(
        OR4_78_Y), .Y(OR4_41_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C2 (.A_DOUT({
        nc19874, nc19875, nc19876, nc19877, nc19878, nc19879, nc19880, 
        nc19881, nc19882, nc19883, nc19884, nc19885, nc19886, nc19887, 
        nc19888, nc19889, nc19890, nc19891, \R_DATA_TEMPR19[5] , 
        \R_DATA_TEMPR19[4] }), .B_DOUT({nc19892, nc19893, nc19894, 
        nc19895, nc19896, nc19897, nc19898, nc19899, nc19900, nc19901, 
        nc19902, nc19903, nc19904, nc19905, nc19906, nc19907, nc19908, 
        nc19909, nc19910, nc19911}), .DB_DETECT(\DB_DETECT[19][2] ), 
        .SB_CORRECT(\SB_CORRECT[19][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C12 (.A_DOUT({
        nc19912, nc19913, nc19914, nc19915, nc19916, nc19917, nc19918, 
        nc19919, nc19920, nc19921, nc19922, nc19923, nc19924, nc19925, 
        nc19926, nc19927, nc19928, nc19929, \R_DATA_TEMPR2[25] , 
        \R_DATA_TEMPR2[24] }), .B_DOUT({nc19930, nc19931, nc19932, 
        nc19933, nc19934, nc19935, nc19936, nc19937, nc19938, nc19939, 
        nc19940, nc19941, nc19942, nc19943, nc19944, nc19945, nc19946, 
        nc19947, nc19948, nc19949}), .DB_DETECT(\DB_DETECT[2][12] ), 
        .SB_CORRECT(\SB_CORRECT[2][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C4 (.A_DOUT({
        nc19950, nc19951, nc19952, nc19953, nc19954, nc19955, nc19956, 
        nc19957, nc19958, nc19959, nc19960, nc19961, nc19962, nc19963, 
        nc19964, nc19965, nc19966, nc19967, \R_DATA_TEMPR29[9] , 
        \R_DATA_TEMPR29[8] }), .B_DOUT({nc19968, nc19969, nc19970, 
        nc19971, nc19972, nc19973, nc19974, nc19975, nc19976, nc19977, 
        nc19978, nc19979, nc19980, nc19981, nc19982, nc19983, nc19984, 
        nc19985, nc19986, nc19987}), .DB_DETECT(\DB_DETECT[29][4] ), 
        .SB_CORRECT(\SB_CORRECT[29][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C18 (.A_DOUT({
        nc19988, nc19989, nc19990, nc19991, nc19992, nc19993, nc19994, 
        nc19995, nc19996, nc19997, nc19998, nc19999, nc20000, nc20001, 
        nc20002, nc20003, nc20004, nc20005, \R_DATA_TEMPR23[37] , 
        \R_DATA_TEMPR23[36] }), .B_DOUT({nc20006, nc20007, nc20008, 
        nc20009, nc20010, nc20011, nc20012, nc20013, nc20014, nc20015, 
        nc20016, nc20017, nc20018, nc20019, nc20020, nc20021, nc20022, 
        nc20023, nc20024, nc20025}), .DB_DETECT(\DB_DETECT[23][18] ), 
        .SB_CORRECT(\SB_CORRECT[23][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_52 (.A(\R_DATA_TEMPR16[21] ), .B(\R_DATA_TEMPR17[21] ), .C(
        \R_DATA_TEMPR18[21] ), .D(\R_DATA_TEMPR19[21] ), .Y(OR4_52_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C16 (.A_DOUT({
        nc20026, nc20027, nc20028, nc20029, nc20030, nc20031, nc20032, 
        nc20033, nc20034, nc20035, nc20036, nc20037, nc20038, nc20039, 
        nc20040, nc20041, nc20042, nc20043, \R_DATA_TEMPR31[33] , 
        \R_DATA_TEMPR31[32] }), .B_DOUT({nc20044, nc20045, nc20046, 
        nc20047, nc20048, nc20049, nc20050, nc20051, nc20052, nc20053, 
        nc20054, nc20055, nc20056, nc20057, nc20058, nc20059, nc20060, 
        nc20061, nc20062, nc20063}), .DB_DETECT(\DB_DETECT[31][16] ), 
        .SB_CORRECT(\SB_CORRECT[31][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_346 (.A(OR4_92_Y), .B(OR2_15_Y), .C(\R_DATA_TEMPR22[11] ), 
        .D(\R_DATA_TEMPR23[11] ), .Y(OR4_346_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C14 (.A_DOUT({
        nc20064, nc20065, nc20066, nc20067, nc20068, nc20069, nc20070, 
        nc20071, nc20072, nc20073, nc20074, nc20075, nc20076, nc20077, 
        nc20078, nc20079, nc20080, nc20081, \R_DATA_TEMPR14[29] , 
        \R_DATA_TEMPR14[28] }), .B_DOUT({nc20082, nc20083, nc20084, 
        nc20085, nc20086, nc20087, nc20088, nc20089, nc20090, nc20091, 
        nc20092, nc20093, nc20094, nc20095, nc20096, nc20097, nc20098, 
        nc20099, nc20100, nc20101}), .DB_DETECT(\DB_DETECT[14][14] ), 
        .SB_CORRECT(\SB_CORRECT[14][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_136 (.A(\R_DATA_TEMPR12[15] ), .B(\R_DATA_TEMPR13[15] ), 
        .C(\R_DATA_TEMPR14[15] ), .D(\R_DATA_TEMPR15[15] ), .Y(
        OR4_136_Y));
    OR2 OR2_20 (.A(\R_DATA_TEMPR20[20] ), .B(\R_DATA_TEMPR21[20] ), .Y(
        OR2_20_Y));
    INV \INVBLKX1[0]  (.A(W_ADDR[14]), .Y(\BLKX1[0] ));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0 (.A_DOUT({nc20102, 
        nc20103, nc20104, nc20105, nc20106, nc20107, nc20108, nc20109, 
        nc20110, nc20111, nc20112, nc20113, nc20114, nc20115, nc20116, 
        nc20117, nc20118, nc20119, \R_DATA_TEMPR1[1] , 
        \R_DATA_TEMPR1[0] }), .B_DOUT({nc20120, nc20121, nc20122, 
        nc20123, nc20124, nc20125, nc20126, nc20127, nc20128, nc20129, 
        nc20130, nc20131, nc20132, nc20133, nc20134, nc20135, nc20136, 
        nc20137, nc20138, nc20139}), .DB_DETECT(\DB_DETECT[1][0] ), 
        .SB_CORRECT(\SB_CORRECT[1][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_16 (.A(\R_DATA_TEMPR20[22] ), .B(\R_DATA_TEMPR21[22] ), .Y(
        OR2_16_Y));
    CFG2 #( .INIT(4'h4) )  CFG2_6 (.A(R_ADDR[16]), .B(R_ADDR[15]), .Y(
        CFG2_6_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C5 (.A_DOUT({nc20140, 
        nc20141, nc20142, nc20143, nc20144, nc20145, nc20146, nc20147, 
        nc20148, nc20149, nc20150, nc20151, nc20152, nc20153, nc20154, 
        nc20155, nc20156, nc20157, \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR5[10] }), .B_DOUT({nc20158, nc20159, nc20160, 
        nc20161, nc20162, nc20163, nc20164, nc20165, nc20166, nc20167, 
        nc20168, nc20169, nc20170, nc20171, nc20172, nc20173, nc20174, 
        nc20175, nc20176, nc20177}), .DB_DETECT(\DB_DETECT[5][5] ), 
        .SB_CORRECT(\SB_CORRECT[5][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C4 (.A_DOUT({nc20178, 
        nc20179, nc20180, nc20181, nc20182, nc20183, nc20184, nc20185, 
        nc20186, nc20187, nc20188, nc20189, nc20190, nc20191, nc20192, 
        nc20193, nc20194, nc20195, \R_DATA_TEMPR8[9] , 
        \R_DATA_TEMPR8[8] }), .B_DOUT({nc20196, nc20197, nc20198, 
        nc20199, nc20200, nc20201, nc20202, nc20203, nc20204, nc20205, 
        nc20206, nc20207, nc20208, nc20209, nc20210, nc20211, nc20212, 
        nc20213, nc20214, nc20215}), .DB_DETECT(\DB_DETECT[8][4] ), 
        .SB_CORRECT(\SB_CORRECT[8][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C19 (.A_DOUT({
        nc20216, nc20217, nc20218, nc20219, nc20220, nc20221, nc20222, 
        nc20223, nc20224, nc20225, nc20226, nc20227, nc20228, nc20229, 
        nc20230, nc20231, nc20232, nc20233, \R_DATA_TEMPR11[39] , 
        \R_DATA_TEMPR11[38] }), .B_DOUT({nc20234, nc20235, nc20236, 
        nc20237, nc20238, nc20239, nc20240, nc20241, nc20242, nc20243, 
        nc20244, nc20245, nc20246, nc20247, nc20248, nc20249, nc20250, 
        nc20251, nc20252, nc20253}), .DB_DETECT(\DB_DETECT[11][19] ), 
        .SB_CORRECT(\SB_CORRECT[11][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C6 (.A_DOUT({
        nc20254, nc20255, nc20256, nc20257, nc20258, nc20259, nc20260, 
        nc20261, nc20262, nc20263, nc20264, nc20265, nc20266, nc20267, 
        nc20268, nc20269, nc20270, nc20271, \R_DATA_TEMPR21[13] , 
        \R_DATA_TEMPR21[12] }), .B_DOUT({nc20272, nc20273, nc20274, 
        nc20275, nc20276, nc20277, nc20278, nc20279, nc20280, nc20281, 
        nc20282, nc20283, nc20284, nc20285, nc20286, nc20287, nc20288, 
        nc20289, nc20290, nc20291}), .DB_DETECT(\DB_DETECT[21][6] ), 
        .SB_CORRECT(\SB_CORRECT[21][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[21][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_27 (.A(\R_DATA_TEMPR20[28] ), .B(\R_DATA_TEMPR21[28] ), .Y(
        OR2_27_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C18 (.A_DOUT({
        nc20292, nc20293, nc20294, nc20295, nc20296, nc20297, nc20298, 
        nc20299, nc20300, nc20301, nc20302, nc20303, nc20304, nc20305, 
        nc20306, nc20307, nc20308, nc20309, \R_DATA_TEMPR3[37] , 
        \R_DATA_TEMPR3[36] }), .B_DOUT({nc20310, nc20311, nc20312, 
        nc20313, nc20314, nc20315, nc20316, nc20317, nc20318, nc20319, 
        nc20320, nc20321, nc20322, nc20323, nc20324, nc20325, nc20326, 
        nc20327, nc20328, nc20329}), .DB_DETECT(\DB_DETECT[3][18] ), 
        .SB_CORRECT(\SB_CORRECT[3][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C14 (.A_DOUT({
        nc20330, nc20331, nc20332, nc20333, nc20334, nc20335, nc20336, 
        nc20337, nc20338, nc20339, nc20340, nc20341, nc20342, nc20343, 
        nc20344, nc20345, nc20346, nc20347, \R_DATA_TEMPR15[29] , 
        \R_DATA_TEMPR15[28] }), .B_DOUT({nc20348, nc20349, nc20350, 
        nc20351, nc20352, nc20353, nc20354, nc20355, nc20356, nc20357, 
        nc20358, nc20359, nc20360, nc20361, nc20362, nc20363, nc20364, 
        nc20365, nc20366, nc20367}), .DB_DETECT(\DB_DETECT[15][14] ), 
        .SB_CORRECT(\SB_CORRECT[15][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[0]  (.A(CFG2_3_Y), .B(
        R_ADDR[17]), .C(R_EN), .Y(\BLKY2[0] ));
    OR4 OR4_203 (.A(\R_DATA_TEMPR24[9] ), .B(\R_DATA_TEMPR25[9] ), .C(
        \R_DATA_TEMPR26[9] ), .D(\R_DATA_TEMPR27[9] ), .Y(OR4_203_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C12 (.A_DOUT({
        nc20368, nc20369, nc20370, nc20371, nc20372, nc20373, nc20374, 
        nc20375, nc20376, nc20377, nc20378, nc20379, nc20380, nc20381, 
        nc20382, nc20383, nc20384, nc20385, \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR7[24] }), .B_DOUT({nc20386, nc20387, nc20388, 
        nc20389, nc20390, nc20391, nc20392, nc20393, nc20394, nc20395, 
        nc20396, nc20397, nc20398, nc20399, nc20400, nc20401, nc20402, 
        nc20403, nc20404, nc20405}), .DB_DETECT(\DB_DETECT[7][12] ), 
        .SB_CORRECT(\SB_CORRECT[7][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_290 (.A(\R_DATA_TEMPR8[25] ), .B(\R_DATA_TEMPR9[25] ), .C(
        \R_DATA_TEMPR10[25] ), .D(\R_DATA_TEMPR11[25] ), .Y(OR4_290_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C6 (.A_DOUT({
        nc20406, nc20407, nc20408, nc20409, nc20410, nc20411, nc20412, 
        nc20413, nc20414, nc20415, nc20416, nc20417, nc20418, nc20419, 
        nc20420, nc20421, nc20422, nc20423, \R_DATA_TEMPR27[13] , 
        \R_DATA_TEMPR27[12] }), .B_DOUT({nc20424, nc20425, nc20426, 
        nc20427, nc20428, nc20429, nc20430, nc20431, nc20432, nc20433, 
        nc20434, nc20435, nc20436, nc20437, nc20438, nc20439, nc20440, 
        nc20441, nc20442, nc20443}), .DB_DETECT(\DB_DETECT[27][6] ), 
        .SB_CORRECT(\SB_CORRECT[27][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_338 (.A(\R_DATA_TEMPR24[29] ), .B(\R_DATA_TEMPR25[29] ), 
        .C(\R_DATA_TEMPR26[29] ), .D(\R_DATA_TEMPR27[29] ), .Y(
        OR4_338_Y));
    OR4 OR4_273 (.A(\R_DATA_TEMPR12[24] ), .B(\R_DATA_TEMPR13[24] ), 
        .C(\R_DATA_TEMPR14[24] ), .D(\R_DATA_TEMPR15[24] ), .Y(
        OR4_273_Y));
    OR4 OR4_322 (.A(\R_DATA_TEMPR12[19] ), .B(\R_DATA_TEMPR13[19] ), 
        .C(\R_DATA_TEMPR14[19] ), .D(\R_DATA_TEMPR15[19] ), .Y(
        OR4_322_Y));
    OR4 OR4_313 (.A(\R_DATA_TEMPR16[25] ), .B(\R_DATA_TEMPR17[25] ), 
        .C(\R_DATA_TEMPR18[25] ), .D(\R_DATA_TEMPR19[25] ), .Y(
        OR4_313_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C19 (.A_DOUT({
        nc20444, nc20445, nc20446, nc20447, nc20448, nc20449, nc20450, 
        nc20451, nc20452, nc20453, nc20454, nc20455, nc20456, nc20457, 
        nc20458, nc20459, nc20460, nc20461, \R_DATA_TEMPR20[39] , 
        \R_DATA_TEMPR20[38] }), .B_DOUT({nc20462, nc20463, nc20464, 
        nc20465, nc20466, nc20467, nc20468, nc20469, nc20470, nc20471, 
        nc20472, nc20473, nc20474, nc20475, nc20476, nc20477, nc20478, 
        nc20479, nc20480, nc20481}), .DB_DETECT(\DB_DETECT[20][19] ), 
        .SB_CORRECT(\SB_CORRECT[20][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_12 (.A(\R_DATA_TEMPR28[17] ), .B(\R_DATA_TEMPR29[17] ), .C(
        \R_DATA_TEMPR30[17] ), .D(\R_DATA_TEMPR31[17] ), .Y(OR4_12_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C11 (.A_DOUT({
        nc20482, nc20483, nc20484, nc20485, nc20486, nc20487, nc20488, 
        nc20489, nc20490, nc20491, nc20492, nc20493, nc20494, nc20495, 
        nc20496, nc20497, nc20498, nc20499, \R_DATA_TEMPR4[23] , 
        \R_DATA_TEMPR4[22] }), .B_DOUT({nc20500, nc20501, nc20502, 
        nc20503, nc20504, nc20505, nc20506, nc20507, nc20508, nc20509, 
        nc20510, nc20511, nc20512, nc20513, nc20514, nc20515, nc20516, 
        nc20517, nc20518, nc20519}), .DB_DETECT(\DB_DETECT[4][11] ), 
        .SB_CORRECT(\SB_CORRECT[4][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_296 (.A(\R_DATA_TEMPR0[22] ), .B(\R_DATA_TEMPR1[22] ), .C(
        \R_DATA_TEMPR2[22] ), .D(\R_DATA_TEMPR3[22] ), .Y(OR4_296_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C12 (.A_DOUT({
        nc20520, nc20521, nc20522, nc20523, nc20524, nc20525, nc20526, 
        nc20527, nc20528, nc20529, nc20530, nc20531, nc20532, nc20533, 
        nc20534, nc20535, nc20536, nc20537, \R_DATA_TEMPR23[25] , 
        \R_DATA_TEMPR23[24] }), .B_DOUT({nc20538, nc20539, nc20540, 
        nc20541, nc20542, nc20543, nc20544, nc20545, nc20546, nc20547, 
        nc20548, nc20549, nc20550, nc20551, nc20552, nc20553, nc20554, 
        nc20555, nc20556, nc20557}), .DB_DETECT(\DB_DETECT[23][12] ), 
        .SB_CORRECT(\SB_CORRECT[23][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_251 (.A(OR4_69_Y), .B(OR2_8_Y), .C(\R_DATA_TEMPR22[6] ), 
        .D(\R_DATA_TEMPR23[6] ), .Y(OR4_251_Y));
    OR4 OR4_79 (.A(\R_DATA_TEMPR24[23] ), .B(\R_DATA_TEMPR25[23] ), .C(
        \R_DATA_TEMPR26[23] ), .D(\R_DATA_TEMPR27[23] ), .Y(OR4_79_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C2 (.A_DOUT({
        nc20558, nc20559, nc20560, nc20561, nc20562, nc20563, nc20564, 
        nc20565, nc20566, nc20567, nc20568, nc20569, nc20570, nc20571, 
        nc20572, nc20573, nc20574, nc20575, \R_DATA_TEMPR13[5] , 
        \R_DATA_TEMPR13[4] }), .B_DOUT({nc20576, nc20577, nc20578, 
        nc20579, nc20580, nc20581, nc20582, nc20583, nc20584, nc20585, 
        nc20586, nc20587, nc20588, nc20589, nc20590, nc20591, nc20592, 
        nc20593, nc20594, nc20595}), .DB_DETECT(\DB_DETECT[13][2] ), 
        .SB_CORRECT(\SB_CORRECT[13][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C10 (.A_DOUT({
        nc20596, nc20597, nc20598, nc20599, nc20600, nc20601, nc20602, 
        nc20603, nc20604, nc20605, nc20606, nc20607, nc20608, nc20609, 
        nc20610, nc20611, nc20612, nc20613, \R_DATA_TEMPR23[21] , 
        \R_DATA_TEMPR23[20] }), .B_DOUT({nc20614, nc20615, nc20616, 
        nc20617, nc20618, nc20619, nc20620, nc20621, nc20622, nc20623, 
        nc20624, nc20625, nc20626, nc20627, nc20628, nc20629, nc20630, 
        nc20631, nc20632, nc20633}), .DB_DETECT(\DB_DETECT[23][10] ), 
        .SB_CORRECT(\SB_CORRECT[23][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_139 (.A(\R_DATA_TEMPR16[3] ), .B(\R_DATA_TEMPR17[3] ), .C(
        \R_DATA_TEMPR18[3] ), .D(\R_DATA_TEMPR19[3] ), .Y(OR4_139_Y));
    OR4 OR4_116 (.A(\R_DATA_TEMPR0[9] ), .B(\R_DATA_TEMPR1[9] ), .C(
        \R_DATA_TEMPR2[9] ), .D(\R_DATA_TEMPR3[9] ), .Y(OR4_116_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C14 (.A_DOUT({
        nc20634, nc20635, nc20636, nc20637, nc20638, nc20639, nc20640, 
        nc20641, nc20642, nc20643, nc20644, nc20645, nc20646, nc20647, 
        nc20648, nc20649, nc20650, nc20651, \R_DATA_TEMPR0[29] , 
        \R_DATA_TEMPR0[28] }), .B_DOUT({nc20652, nc20653, nc20654, 
        nc20655, nc20656, nc20657, nc20658, nc20659, nc20660, nc20661, 
        nc20662, nc20663, nc20664, nc20665, nc20666, nc20667, nc20668, 
        nc20669, nc20670, nc20671}), .DB_DETECT(\DB_DETECT[0][14] ), 
        .SB_CORRECT(\SB_CORRECT[0][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_144 (.A(\R_DATA_TEMPR16[30] ), .B(\R_DATA_TEMPR17[30] ), 
        .C(\R_DATA_TEMPR18[30] ), .D(\R_DATA_TEMPR19[30] ), .Y(
        OR4_144_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C3 (.A_DOUT({
        nc20672, nc20673, nc20674, nc20675, nc20676, nc20677, nc20678, 
        nc20679, nc20680, nc20681, nc20682, nc20683, nc20684, nc20685, 
        nc20686, nc20687, nc20688, nc20689, \R_DATA_TEMPR28[7] , 
        \R_DATA_TEMPR28[6] }), .B_DOUT({nc20690, nc20691, nc20692, 
        nc20693, nc20694, nc20695, nc20696, nc20697, nc20698, nc20699, 
        nc20700, nc20701, nc20702, nc20703, nc20704, nc20705, nc20706, 
        nc20707, nc20708, nc20709}), .DB_DETECT(\DB_DETECT[28][3] ), 
        .SB_CORRECT(\SB_CORRECT[28][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[28][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C4 (.A_DOUT({
        nc20710, nc20711, nc20712, nc20713, nc20714, nc20715, nc20716, 
        nc20717, nc20718, nc20719, nc20720, nc20721, nc20722, nc20723, 
        nc20724, nc20725, nc20726, nc20727, \R_DATA_TEMPR15[9] , 
        \R_DATA_TEMPR15[8] }), .B_DOUT({nc20728, nc20729, nc20730, 
        nc20731, nc20732, nc20733, nc20734, nc20735, nc20736, nc20737, 
        nc20738, nc20739, nc20740, nc20741, nc20742, nc20743, nc20744, 
        nc20745, nc20746, nc20747}), .DB_DETECT(\DB_DETECT[15][4] ), 
        .SB_CORRECT(\SB_CORRECT[15][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C17 (.A_DOUT({
        nc20748, nc20749, nc20750, nc20751, nc20752, nc20753, nc20754, 
        nc20755, nc20756, nc20757, nc20758, nc20759, nc20760, nc20761, 
        nc20762, nc20763, nc20764, nc20765, \R_DATA_TEMPR16[35] , 
        \R_DATA_TEMPR16[34] }), .B_DOUT({nc20766, nc20767, nc20768, 
        nc20769, nc20770, nc20771, nc20772, nc20773, nc20774, nc20775, 
        nc20776, nc20777, nc20778, nc20779, nc20780, nc20781, nc20782, 
        nc20783, nc20784, nc20785}), .DB_DETECT(\DB_DETECT[16][17] ), 
        .SB_CORRECT(\SB_CORRECT[16][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C12 (.A_DOUT({
        nc20786, nc20787, nc20788, nc20789, nc20790, nc20791, nc20792, 
        nc20793, nc20794, nc20795, nc20796, nc20797, nc20798, nc20799, 
        nc20800, nc20801, nc20802, nc20803, \R_DATA_TEMPR5[25] , 
        \R_DATA_TEMPR5[24] }), .B_DOUT({nc20804, nc20805, nc20806, 
        nc20807, nc20808, nc20809, nc20810, nc20811, nc20812, nc20813, 
        nc20814, nc20815, nc20816, nc20817, nc20818, nc20819, nc20820, 
        nc20821, nc20822, nc20823}), .DB_DETECT(\DB_DETECT[5][12] ), 
        .SB_CORRECT(\SB_CORRECT[5][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[32]  (.A(OR4_345_Y), .B(OR4_330_Y), .C(OR4_282_Y), 
        .D(OR4_124_Y), .Y(R_DATA[32]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C16 (.A_DOUT({
        nc20824, nc20825, nc20826, nc20827, nc20828, nc20829, nc20830, 
        nc20831, nc20832, nc20833, nc20834, nc20835, nc20836, nc20837, 
        nc20838, nc20839, nc20840, nc20841, \R_DATA_TEMPR13[33] , 
        \R_DATA_TEMPR13[32] }), .B_DOUT({nc20842, nc20843, nc20844, 
        nc20845, nc20846, nc20847, nc20848, nc20849, nc20850, nc20851, 
        nc20852, nc20853, nc20854, nc20855, nc20856, nc20857, nc20858, 
        nc20859, nc20860, nc20861}), .DB_DETECT(\DB_DETECT[13][16] ), 
        .SB_CORRECT(\SB_CORRECT[13][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C1 (.A_DOUT({
        nc20862, nc20863, nc20864, nc20865, nc20866, nc20867, nc20868, 
        nc20869, nc20870, nc20871, nc20872, nc20873, nc20874, nc20875, 
        nc20876, nc20877, nc20878, nc20879, \R_DATA_TEMPR21[3] , 
        \R_DATA_TEMPR21[2] }), .B_DOUT({nc20880, nc20881, nc20882, 
        nc20883, nc20884, nc20885, nc20886, nc20887, nc20888, nc20889, 
        nc20890, nc20891, nc20892, nc20893, nc20894, nc20895, nc20896, 
        nc20897, nc20898, nc20899}), .DB_DETECT(\DB_DETECT[21][1] ), 
        .SB_CORRECT(\SB_CORRECT[21][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[21][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C10 (.A_DOUT({
        nc20900, nc20901, nc20902, nc20903, nc20904, nc20905, nc20906, 
        nc20907, nc20908, nc20909, nc20910, nc20911, nc20912, nc20913, 
        nc20914, nc20915, nc20916, nc20917, \R_DATA_TEMPR19[21] , 
        \R_DATA_TEMPR19[20] }), .B_DOUT({nc20918, nc20919, nc20920, 
        nc20921, nc20922, nc20923, nc20924, nc20925, nc20926, nc20927, 
        nc20928, nc20929, nc20930, nc20931, nc20932, nc20933, nc20934, 
        nc20935, nc20936, nc20937}), .DB_DETECT(\DB_DETECT[19][10] ), 
        .SB_CORRECT(\SB_CORRECT[19][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_220 (.A(\R_DATA_TEMPR24[0] ), .B(\R_DATA_TEMPR25[0] ), .C(
        \R_DATA_TEMPR26[0] ), .D(\R_DATA_TEMPR27[0] ), .Y(OR4_220_Y));
    OR4 OR4_318 (.A(\R_DATA_TEMPR12[16] ), .B(\R_DATA_TEMPR13[16] ), 
        .C(\R_DATA_TEMPR14[16] ), .D(\R_DATA_TEMPR15[16] ), .Y(
        OR4_318_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C15 (.A_DOUT({
        nc20938, nc20939, nc20940, nc20941, nc20942, nc20943, nc20944, 
        nc20945, nc20946, nc20947, nc20948, nc20949, nc20950, nc20951, 
        nc20952, nc20953, nc20954, nc20955, \R_DATA_TEMPR19[31] , 
        \R_DATA_TEMPR19[30] }), .B_DOUT({nc20956, nc20957, nc20958, 
        nc20959, nc20960, nc20961, nc20962, nc20963, nc20964, nc20965, 
        nc20966, nc20967, nc20968, nc20969, nc20970, nc20971, nc20972, 
        nc20973, nc20974, nc20975}), .DB_DETECT(\DB_DETECT[19][15] ), 
        .SB_CORRECT(\SB_CORRECT[19][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C8 (.A_DOUT({
        nc20976, nc20977, nc20978, nc20979, nc20980, nc20981, nc20982, 
        nc20983, nc20984, nc20985, nc20986, nc20987, nc20988, nc20989, 
        nc20990, nc20991, nc20992, nc20993, \R_DATA_TEMPR20[17] , 
        \R_DATA_TEMPR20[16] }), .B_DOUT({nc20994, nc20995, nc20996, 
        nc20997, nc20998, nc20999, nc21000, nc21001, nc21002, nc21003, 
        nc21004, nc21005, nc21006, nc21007, nc21008, nc21009, nc21010, 
        nc21011, nc21012, nc21013}), .DB_DETECT(\DB_DETECT[20][8] ), 
        .SB_CORRECT(\SB_CORRECT[20][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_10 (.A(\R_DATA_TEMPR20[23] ), .B(\R_DATA_TEMPR21[23] ), .Y(
        OR2_10_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C18 (.A_DOUT({
        nc21014, nc21015, nc21016, nc21017, nc21018, nc21019, nc21020, 
        nc21021, nc21022, nc21023, nc21024, nc21025, nc21026, nc21027, 
        nc21028, nc21029, nc21030, nc21031, \R_DATA_TEMPR20[37] , 
        \R_DATA_TEMPR20[36] }), .B_DOUT({nc21032, nc21033, nc21034, 
        nc21035, nc21036, nc21037, nc21038, nc21039, nc21040, nc21041, 
        nc21042, nc21043, nc21044, nc21045, nc21046, nc21047, nc21048, 
        nc21049, nc21050, nc21051}), .DB_DETECT(\DB_DETECT[20][18] ), 
        .SB_CORRECT(\SB_CORRECT[20][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[3]  (.A(OR4_89_Y), .B(OR4_180_Y), .C(OR4_151_Y), 
        .D(OR4_179_Y), .Y(R_DATA[3]));
    OR2 OR2_17 (.A(\R_DATA_TEMPR20[34] ), .B(\R_DATA_TEMPR21[34] ), .Y(
        OR2_17_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0 (.A_DOUT({
        nc21052, nc21053, nc21054, nc21055, nc21056, nc21057, nc21058, 
        nc21059, nc21060, nc21061, nc21062, nc21063, nc21064, nc21065, 
        nc21066, nc21067, nc21068, nc21069, \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR15[0] }), .B_DOUT({nc21070, nc21071, nc21072, 
        nc21073, nc21074, nc21075, nc21076, nc21077, nc21078, nc21079, 
        nc21080, nc21081, nc21082, nc21083, nc21084, nc21085, nc21086, 
        nc21087, nc21088, nc21089}), .DB_DETECT(\DB_DETECT[15][0] ), 
        .SB_CORRECT(\SB_CORRECT[15][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C2 (.A_DOUT({nc21090, 
        nc21091, nc21092, nc21093, nc21094, nc21095, nc21096, nc21097, 
        nc21098, nc21099, nc21100, nc21101, nc21102, nc21103, nc21104, 
        nc21105, nc21106, nc21107, \R_DATA_TEMPR2[5] , 
        \R_DATA_TEMPR2[4] }), .B_DOUT({nc21108, nc21109, nc21110, 
        nc21111, nc21112, nc21113, nc21114, nc21115, nc21116, nc21117, 
        nc21118, nc21119, nc21120, nc21121, nc21122, nc21123, nc21124, 
        nc21125, nc21126, nc21127}), .DB_DETECT(\DB_DETECT[2][2] ), 
        .SB_CORRECT(\SB_CORRECT[2][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C11 (.A_DOUT({
        nc21128, nc21129, nc21130, nc21131, nc21132, nc21133, nc21134, 
        nc21135, nc21136, nc21137, nc21138, nc21139, nc21140, nc21141, 
        nc21142, nc21143, nc21144, nc21145, \R_DATA_TEMPR18[23] , 
        \R_DATA_TEMPR18[22] }), .B_DOUT({nc21146, nc21147, nc21148, 
        nc21149, nc21150, nc21151, nc21152, nc21153, nc21154, nc21155, 
        nc21156, nc21157, nc21158, nc21159, nc21160, nc21161, nc21162, 
        nc21163, nc21164, nc21165}), .DB_DETECT(\DB_DETECT[18][11] ), 
        .SB_CORRECT(\SB_CORRECT[18][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C19 (.A_DOUT({
        nc21166, nc21167, nc21168, nc21169, nc21170, nc21171, nc21172, 
        nc21173, nc21174, nc21175, nc21176, nc21177, nc21178, nc21179, 
        nc21180, nc21181, nc21182, nc21183, \R_DATA_TEMPR24[39] , 
        \R_DATA_TEMPR24[38] }), .B_DOUT({nc21184, nc21185, nc21186, 
        nc21187, nc21188, nc21189, nc21190, nc21191, nc21192, nc21193, 
        nc21194, nc21195, nc21196, nc21197, nc21198, nc21199, nc21200, 
        nc21201, nc21202, nc21203}), .DB_DETECT(\DB_DETECT[24][19] ), 
        .SB_CORRECT(\SB_CORRECT[24][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C4 (.A_DOUT({
        nc21204, nc21205, nc21206, nc21207, nc21208, nc21209, nc21210, 
        nc21211, nc21212, nc21213, nc21214, nc21215, nc21216, nc21217, 
        nc21218, nc21219, nc21220, nc21221, \R_DATA_TEMPR24[9] , 
        \R_DATA_TEMPR24[8] }), .B_DOUT({nc21222, nc21223, nc21224, 
        nc21225, nc21226, nc21227, nc21228, nc21229, nc21230, nc21231, 
        nc21232, nc21233, nc21234, nc21235, nc21236, nc21237, nc21238, 
        nc21239, nc21240, nc21241}), .DB_DETECT(\DB_DETECT[24][4] ), 
        .SB_CORRECT(\SB_CORRECT[24][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_226 (.A(\R_DATA_TEMPR12[4] ), .B(\R_DATA_TEMPR13[4] ), .C(
        \R_DATA_TEMPR14[4] ), .D(\R_DATA_TEMPR15[4] ), .Y(OR4_226_Y));
    OR4 OR4_119 (.A(\R_DATA_TEMPR24[34] ), .B(\R_DATA_TEMPR25[34] ), 
        .C(\R_DATA_TEMPR26[34] ), .D(\R_DATA_TEMPR27[34] ), .Y(
        OR4_119_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C8 (.A_DOUT({
        nc21242, nc21243, nc21244, nc21245, nc21246, nc21247, nc21248, 
        nc21249, nc21250, nc21251, nc21252, nc21253, nc21254, nc21255, 
        nc21256, nc21257, nc21258, nc21259, \R_DATA_TEMPR27[17] , 
        \R_DATA_TEMPR27[16] }), .B_DOUT({nc21260, nc21261, nc21262, 
        nc21263, nc21264, nc21265, nc21266, nc21267, nc21268, nc21269, 
        nc21270, nc21271, nc21272, nc21273, nc21274, nc21275, nc21276, 
        nc21277, nc21278, nc21279}), .DB_DETECT(\DB_DETECT[27][8] ), 
        .SB_CORRECT(\SB_CORRECT[27][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C8 (.A_DOUT({
        nc21280, nc21281, nc21282, nc21283, nc21284, nc21285, nc21286, 
        nc21287, nc21288, nc21289, nc21290, nc21291, nc21292, nc21293, 
        nc21294, nc21295, nc21296, nc21297, \R_DATA_TEMPR19[17] , 
        \R_DATA_TEMPR19[16] }), .B_DOUT({nc21298, nc21299, nc21300, 
        nc21301, nc21302, nc21303, nc21304, nc21305, nc21306, nc21307, 
        nc21308, nc21309, nc21310, nc21311, nc21312, nc21313, nc21314, 
        nc21315, nc21316, nc21317}), .DB_DETECT(\DB_DETECT[19][8] ), 
        .SB_CORRECT(\SB_CORRECT[19][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[19][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_72 (.A(\R_DATA_TEMPR12[12] ), .B(\R_DATA_TEMPR13[12] ), .C(
        \R_DATA_TEMPR14[12] ), .D(\R_DATA_TEMPR15[12] ), .Y(OR4_72_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C19 (.A_DOUT({
        nc21318, nc21319, nc21320, nc21321, nc21322, nc21323, nc21324, 
        nc21325, nc21326, nc21327, nc21328, nc21329, nc21330, nc21331, 
        nc21332, nc21333, nc21334, nc21335, \R_DATA_TEMPR25[39] , 
        \R_DATA_TEMPR25[38] }), .B_DOUT({nc21336, nc21337, nc21338, 
        nc21339, nc21340, nc21341, nc21342, nc21343, nc21344, nc21345, 
        nc21346, nc21347, nc21348, nc21349, nc21350, nc21351, nc21352, 
        nc21353, nc21354, nc21355}), .DB_DETECT(\DB_DETECT[25][19] ), 
        .SB_CORRECT(\SB_CORRECT[25][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C19 (.A_DOUT({
        nc21356, nc21357, nc21358, nc21359, nc21360, nc21361, nc21362, 
        nc21363, nc21364, nc21365, nc21366, nc21367, nc21368, nc21369, 
        nc21370, nc21371, nc21372, nc21373, \R_DATA_TEMPR2[39] , 
        \R_DATA_TEMPR2[38] }), .B_DOUT({nc21374, nc21375, nc21376, 
        nc21377, nc21378, nc21379, nc21380, nc21381, nc21382, nc21383, 
        nc21384, nc21385, nc21386, nc21387, nc21388, nc21389, nc21390, 
        nc21391, nc21392, nc21393}), .DB_DETECT(\DB_DETECT[2][19] ), 
        .SB_CORRECT(\SB_CORRECT[2][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C2 (.A_DOUT({nc21394, 
        nc21395, nc21396, nc21397, nc21398, nc21399, nc21400, nc21401, 
        nc21402, nc21403, nc21404, nc21405, nc21406, nc21407, nc21408, 
        nc21409, nc21410, nc21411, \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR7[4] }), .B_DOUT({nc21412, nc21413, nc21414, 
        nc21415, nc21416, nc21417, nc21418, nc21419, nc21420, nc21421, 
        nc21422, nc21423, nc21424, nc21425, nc21426, nc21427, nc21428, 
        nc21429, nc21430, nc21431}), .DB_DETECT(\DB_DETECT[7][2] ), 
        .SB_CORRECT(\SB_CORRECT[7][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C8 (.A_DOUT({nc21432, 
        nc21433, nc21434, nc21435, nc21436, nc21437, nc21438, nc21439, 
        nc21440, nc21441, nc21442, nc21443, nc21444, nc21445, nc21446, 
        nc21447, nc21448, nc21449, \R_DATA_TEMPR3[17] , 
        \R_DATA_TEMPR3[16] }), .B_DOUT({nc21450, nc21451, nc21452, 
        nc21453, nc21454, nc21455, nc21456, nc21457, nc21458, nc21459, 
        nc21460, nc21461, nc21462, nc21463, nc21464, nc21465, nc21466, 
        nc21467, nc21468, nc21469}), .DB_DETECT(\DB_DETECT[3][8] ), 
        .SB_CORRECT(\SB_CORRECT[3][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_351 (.A(OR4_32_Y), .B(OR2_20_Y), .C(\R_DATA_TEMPR22[20] ), 
        .D(\R_DATA_TEMPR23[20] ), .Y(OR4_351_Y));
    OR2 OR2_28 (.A(\R_DATA_TEMPR20[19] ), .B(\R_DATA_TEMPR21[19] ), .Y(
        OR2_28_Y));
    OR4 \OR4_R_DATA[33]  (.A(OR4_301_Y), .B(OR4_205_Y), .C(OR4_191_Y), 
        .D(OR4_176_Y), .Y(R_DATA[33]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C4 (.A_DOUT({
        nc21470, nc21471, nc21472, nc21473, nc21474, nc21475, nc21476, 
        nc21477, nc21478, nc21479, nc21480, nc21481, nc21482, nc21483, 
        nc21484, nc21485, nc21486, nc21487, \R_DATA_TEMPR12[9] , 
        \R_DATA_TEMPR12[8] }), .B_DOUT({nc21488, nc21489, nc21490, 
        nc21491, nc21492, nc21493, nc21494, nc21495, nc21496, nc21497, 
        nc21498, nc21499, nc21500, nc21501, nc21502, nc21503, nc21504, 
        nc21505, nc21506, nc21507}), .DB_DETECT(\DB_DETECT[12][4] ), 
        .SB_CORRECT(\SB_CORRECT[12][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C2 (.A_DOUT({
        nc21508, nc21509, nc21510, nc21511, nc21512, nc21513, nc21514, 
        nc21515, nc21516, nc21517, nc21518, nc21519, nc21520, nc21521, 
        nc21522, nc21523, nc21524, nc21525, \R_DATA_TEMPR12[5] , 
        \R_DATA_TEMPR12[4] }), .B_DOUT({nc21526, nc21527, nc21528, 
        nc21529, nc21530, nc21531, nc21532, nc21533, nc21534, nc21535, 
        nc21536, nc21537, nc21538, nc21539, nc21540, nc21541, nc21542, 
        nc21543, nc21544, nc21545}), .DB_DETECT(\DB_DETECT[12][2] ), 
        .SB_CORRECT(\SB_CORRECT[12][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C13 (.A_DOUT({
        nc21546, nc21547, nc21548, nc21549, nc21550, nc21551, nc21552, 
        nc21553, nc21554, nc21555, nc21556, nc21557, nc21558, nc21559, 
        nc21560, nc21561, nc21562, nc21563, \R_DATA_TEMPR13[27] , 
        \R_DATA_TEMPR13[26] }), .B_DOUT({nc21564, nc21565, nc21566, 
        nc21567, nc21568, nc21569, nc21570, nc21571, nc21572, nc21573, 
        nc21574, nc21575, nc21576, nc21577, nc21578, nc21579, nc21580, 
        nc21581, nc21582, nc21583}), .DB_DETECT(\DB_DETECT[13][13] ), 
        .SB_CORRECT(\SB_CORRECT[13][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[13][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C6 (.A_DOUT({
        nc21584, nc21585, nc21586, nc21587, nc21588, nc21589, nc21590, 
        nc21591, nc21592, nc21593, nc21594, nc21595, nc21596, nc21597, 
        nc21598, nc21599, nc21600, nc21601, \R_DATA_TEMPR24[13] , 
        \R_DATA_TEMPR24[12] }), .B_DOUT({nc21602, nc21603, nc21604, 
        nc21605, nc21606, nc21607, nc21608, nc21609, nc21610, nc21611, 
        nc21612, nc21613, nc21614, nc21615, nc21616, nc21617, nc21618, 
        nc21619, nc21620, nc21621}), .DB_DETECT(\DB_DETECT[24][6] ), 
        .SB_CORRECT(\SB_CORRECT[24][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[25]  (.A(OR4_285_Y), .B(OR4_97_Y), .C(OR4_230_Y), 
        .D(OR4_133_Y), .Y(R_DATA[25]));
    OR4 OR4_283 (.A(\R_DATA_TEMPR4[0] ), .B(\R_DATA_TEMPR5[0] ), .C(
        \R_DATA_TEMPR6[0] ), .D(\R_DATA_TEMPR7[0] ), .Y(OR4_283_Y));
    OR4 OR4_96 (.A(\R_DATA_TEMPR0[15] ), .B(\R_DATA_TEMPR1[15] ), .C(
        \R_DATA_TEMPR2[15] ), .D(\R_DATA_TEMPR3[15] ), .Y(OR4_96_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C5 (.A_DOUT({
        nc21622, nc21623, nc21624, nc21625, nc21626, nc21627, nc21628, 
        nc21629, nc21630, nc21631, nc21632, nc21633, nc21634, nc21635, 
        nc21636, nc21637, nc21638, nc21639, \R_DATA_TEMPR29[11] , 
        \R_DATA_TEMPR29[10] }), .B_DOUT({nc21640, nc21641, nc21642, 
        nc21643, nc21644, nc21645, nc21646, nc21647, nc21648, nc21649, 
        nc21650, nc21651, nc21652, nc21653, nc21654, nc21655, nc21656, 
        nc21657, nc21658, nc21659}), .DB_DETECT(\DB_DETECT[29][5] ), 
        .SB_CORRECT(\SB_CORRECT[29][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[29][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C12 (.A_DOUT({
        nc21660, nc21661, nc21662, nc21663, nc21664, nc21665, nc21666, 
        nc21667, nc21668, nc21669, nc21670, nc21671, nc21672, nc21673, 
        nc21674, nc21675, nc21676, nc21677, \R_DATA_TEMPR20[25] , 
        \R_DATA_TEMPR20[24] }), .B_DOUT({nc21678, nc21679, nc21680, 
        nc21681, nc21682, nc21683, nc21684, nc21685, nc21686, nc21687, 
        nc21688, nc21689, nc21690, nc21691, nc21692, nc21693, nc21694, 
        nc21695, nc21696, nc21697}), .DB_DETECT(\DB_DETECT[20][12] ), 
        .SB_CORRECT(\SB_CORRECT[20][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C6 (.A_DOUT({nc21698, 
        nc21699, nc21700, nc21701, nc21702, nc21703, nc21704, nc21705, 
        nc21706, nc21707, nc21708, nc21709, nc21710, nc21711, nc21712, 
        nc21713, nc21714, nc21715, \R_DATA_TEMPR2[13] , 
        \R_DATA_TEMPR2[12] }), .B_DOUT({nc21716, nc21717, nc21718, 
        nc21719, nc21720, nc21721, nc21722, nc21723, nc21724, nc21725, 
        nc21726, nc21727, nc21728, nc21729, nc21730, nc21731, nc21732, 
        nc21733, nc21734, nc21735}), .DB_DETECT(\DB_DETECT[2][6] ), 
        .SB_CORRECT(\SB_CORRECT[2][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C10 (.A_DOUT({
        nc21736, nc21737, nc21738, nc21739, nc21740, nc21741, nc21742, 
        nc21743, nc21744, nc21745, nc21746, nc21747, nc21748, nc21749, 
        nc21750, nc21751, nc21752, nc21753, \R_DATA_TEMPR20[21] , 
        \R_DATA_TEMPR20[20] }), .B_DOUT({nc21754, nc21755, nc21756, 
        nc21757, nc21758, nc21759, nc21760, nc21761, nc21762, nc21763, 
        nc21764, nc21765, nc21766, nc21767, nc21768, nc21769, nc21770, 
        nc21771, nc21772, nc21773}), .DB_DETECT(\DB_DETECT[20][10] ), 
        .SB_CORRECT(\SB_CORRECT[20][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C18 (.A_DOUT({
        nc21774, nc21775, nc21776, nc21777, nc21778, nc21779, nc21780, 
        nc21781, nc21782, nc21783, nc21784, nc21785, nc21786, nc21787, 
        nc21788, nc21789, nc21790, nc21791, \R_DATA_TEMPR24[37] , 
        \R_DATA_TEMPR24[36] }), .B_DOUT({nc21792, nc21793, nc21794, 
        nc21795, nc21796, nc21797, nc21798, nc21799, nc21800, nc21801, 
        nc21802, nc21803, nc21804, nc21805, nc21806, nc21807, nc21808, 
        nc21809, nc21810, nc21811}), .DB_DETECT(\DB_DETECT[24][18] ), 
        .SB_CORRECT(\SB_CORRECT[24][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1 (.A_DOUT({nc21812, 
        nc21813, nc21814, nc21815, nc21816, nc21817, nc21818, nc21819, 
        nc21820, nc21821, nc21822, nc21823, nc21824, nc21825, nc21826, 
        nc21827, nc21828, nc21829, \R_DATA_TEMPR9[3] , 
        \R_DATA_TEMPR9[2] }), .B_DOUT({nc21830, nc21831, nc21832, 
        nc21833, nc21834, nc21835, nc21836, nc21837, nc21838, nc21839, 
        nc21840, nc21841, nc21842, nc21843, nc21844, nc21845, nc21846, 
        nc21847, nc21848, nc21849}), .DB_DETECT(\DB_DETECT[9][1] ), 
        .SB_CORRECT(\SB_CORRECT[9][1] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][1] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[3], W_DATA[2]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[1]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C19 (.A_DOUT({
        nc21850, nc21851, nc21852, nc21853, nc21854, nc21855, nc21856, 
        nc21857, nc21858, nc21859, nc21860, nc21861, nc21862, nc21863, 
        nc21864, nc21865, nc21866, nc21867, \R_DATA_TEMPR7[39] , 
        \R_DATA_TEMPR7[38] }), .B_DOUT({nc21868, nc21869, nc21870, 
        nc21871, nc21872, nc21873, nc21874, nc21875, nc21876, nc21877, 
        nc21878, nc21879, nc21880, nc21881, nc21882, nc21883, nc21884, 
        nc21885, nc21886, nc21887}), .DB_DETECT(\DB_DETECT[7][19] ), 
        .SB_CORRECT(\SB_CORRECT[7][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_54 (.A(\R_DATA_TEMPR0[33] ), .B(\R_DATA_TEMPR1[33] ), .C(
        \R_DATA_TEMPR2[33] ), .D(\R_DATA_TEMPR3[33] ), .Y(OR4_54_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C5 (.A_DOUT({nc21888, 
        nc21889, nc21890, nc21891, nc21892, nc21893, nc21894, nc21895, 
        nc21896, nc21897, nc21898, nc21899, nc21900, nc21901, nc21902, 
        nc21903, nc21904, nc21905, \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR2[10] }), .B_DOUT({nc21906, nc21907, nc21908, 
        nc21909, nc21910, nc21911, nc21912, nc21913, nc21914, nc21915, 
        nc21916, nc21917, nc21918, nc21919, nc21920, nc21921, nc21922, 
        nc21923, nc21924, nc21925}), .DB_DETECT(\DB_DETECT[2][5] ), 
        .SB_CORRECT(\SB_CORRECT[2][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[2][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C18 (.A_DOUT({
        nc21926, nc21927, nc21928, nc21929, nc21930, nc21931, nc21932, 
        nc21933, nc21934, nc21935, nc21936, nc21937, nc21938, nc21939, 
        nc21940, nc21941, nc21942, nc21943, \R_DATA_TEMPR0[37] , 
        \R_DATA_TEMPR0[36] }), .B_DOUT({nc21944, nc21945, nc21946, 
        nc21947, nc21948, nc21949, nc21950, nc21951, nc21952, nc21953, 
        nc21954, nc21955, nc21956, nc21957, nc21958, nc21959, nc21960, 
        nc21961, nc21962, nc21963}), .DB_DETECT(\DB_DETECT[0][18] ), 
        .SB_CORRECT(\SB_CORRECT[0][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_3 (.A(OR4_155_Y), .B(OR2_39_Y), .C(\R_DATA_TEMPR22[29] ), 
        .D(\R_DATA_TEMPR23[29] ), .Y(OR4_3_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C18 (.A_DOUT({
        nc21964, nc21965, nc21966, nc21967, nc21968, nc21969, nc21970, 
        nc21971, nc21972, nc21973, nc21974, nc21975, nc21976, nc21977, 
        nc21978, nc21979, nc21980, nc21981, \R_DATA_TEMPR25[37] , 
        \R_DATA_TEMPR25[36] }), .B_DOUT({nc21982, nc21983, nc21984, 
        nc21985, nc21986, nc21987, nc21988, nc21989, nc21990, nc21991, 
        nc21992, nc21993, nc21994, nc21995, nc21996, nc21997, nc21998, 
        nc21999, nc22000, nc22001}), .DB_DETECT(\DB_DETECT[25][18] ), 
        .SB_CORRECT(\SB_CORRECT[25][18] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][18] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[37], W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[18]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C17 (.A_DOUT({
        nc22002, nc22003, nc22004, nc22005, nc22006, nc22007, nc22008, 
        nc22009, nc22010, nc22011, nc22012, nc22013, nc22014, nc22015, 
        nc22016, nc22017, nc22018, nc22019, \R_DATA_TEMPR23[35] , 
        \R_DATA_TEMPR23[34] }), .B_DOUT({nc22020, nc22021, nc22022, 
        nc22023, nc22024, nc22025, nc22026, nc22027, nc22028, nc22029, 
        nc22030, nc22031, nc22032, nc22033, nc22034, nc22035, nc22036, 
        nc22037, nc22038, nc22039}), .DB_DETECT(\DB_DETECT[23][17] ), 
        .SB_CORRECT(\SB_CORRECT[23][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C8 (.A_DOUT({
        nc22040, nc22041, nc22042, nc22043, nc22044, nc22045, nc22046, 
        nc22047, nc22048, nc22049, nc22050, nc22051, nc22052, nc22053, 
        nc22054, nc22055, nc22056, nc22057, \R_DATA_TEMPR23[17] , 
        \R_DATA_TEMPR23[16] }), .B_DOUT({nc22058, nc22059, nc22060, 
        nc22061, nc22062, nc22063, nc22064, nc22065, nc22066, nc22067, 
        nc22068, nc22069, nc22070, nc22071, nc22072, nc22073, nc22074, 
        nc22075, nc22076, nc22077}), .DB_DETECT(\DB_DETECT[23][8] ), 
        .SB_CORRECT(\SB_CORRECT[23][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C16 (.A_DOUT({
        nc22078, nc22079, nc22080, nc22081, nc22082, nc22083, nc22084, 
        nc22085, nc22086, nc22087, nc22088, nc22089, nc22090, nc22091, 
        nc22092, nc22093, nc22094, nc22095, \R_DATA_TEMPR10[33] , 
        \R_DATA_TEMPR10[32] }), .B_DOUT({nc22096, nc22097, nc22098, 
        nc22099, nc22100, nc22101, nc22102, nc22103, nc22104, nc22105, 
        nc22106, nc22107, nc22108, nc22109, nc22110, nc22111, nc22112, 
        nc22113, nc22114, nc22115}), .DB_DETECT(\DB_DETECT[10][16] ), 
        .SB_CORRECT(\SB_CORRECT[10][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_161 (.A(\R_DATA_TEMPR16[27] ), .B(\R_DATA_TEMPR17[27] ), 
        .C(\R_DATA_TEMPR18[27] ), .D(\R_DATA_TEMPR19[27] ), .Y(
        OR4_161_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C4 (.A_DOUT({
        nc22116, nc22117, nc22118, nc22119, nc22120, nc22121, nc22122, 
        nc22123, nc22124, nc22125, nc22126, nc22127, nc22128, nc22129, 
        nc22130, nc22131, nc22132, nc22133, \R_DATA_TEMPR16[9] , 
        \R_DATA_TEMPR16[8] }), .B_DOUT({nc22134, nc22135, nc22136, 
        nc22137, nc22138, nc22139, nc22140, nc22141, nc22142, nc22143, 
        nc22144, nc22145, nc22146, nc22147, nc22148, nc22149, nc22150, 
        nc22151, nc22152, nc22153}), .DB_DETECT(\DB_DETECT[16][4] ), 
        .SB_CORRECT(\SB_CORRECT[16][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C17 (.A_DOUT({
        nc22154, nc22155, nc22156, nc22157, nc22158, nc22159, nc22160, 
        nc22161, nc22162, nc22163, nc22164, nc22165, nc22166, nc22167, 
        nc22168, nc22169, nc22170, nc22171, \R_DATA_TEMPR9[35] , 
        \R_DATA_TEMPR9[34] }), .B_DOUT({nc22172, nc22173, nc22174, 
        nc22175, nc22176, nc22177, nc22178, nc22179, nc22180, nc22181, 
        nc22182, nc22183, nc22184, nc22185, nc22186, nc22187, nc22188, 
        nc22189, nc22190, nc22191}), .DB_DETECT(\DB_DETECT[9][17] ), 
        .SB_CORRECT(\SB_CORRECT[9][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_237 (.A(\R_DATA_TEMPR28[11] ), .B(\R_DATA_TEMPR29[11] ), 
        .C(\R_DATA_TEMPR30[11] ), .D(\R_DATA_TEMPR31[11] ), .Y(
        OR4_237_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C2 (.A_DOUT({
        nc22192, nc22193, nc22194, nc22195, nc22196, nc22197, nc22198, 
        nc22199, nc22200, nc22201, nc22202, nc22203, nc22204, nc22205, 
        nc22206, nc22207, nc22208, nc22209, \R_DATA_TEMPR10[5] , 
        \R_DATA_TEMPR10[4] }), .B_DOUT({nc22210, nc22211, nc22212, 
        nc22213, nc22214, nc22215, nc22216, nc22217, nc22218, nc22219, 
        nc22220, nc22221, nc22222, nc22223, nc22224, nc22225, nc22226, 
        nc22227, nc22228, nc22229}), .DB_DETECT(\DB_DETECT[10][2] ), 
        .SB_CORRECT(\SB_CORRECT[10][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C17 (.A_DOUT({
        nc22230, nc22231, nc22232, nc22233, nc22234, nc22235, nc22236, 
        nc22237, nc22238, nc22239, nc22240, nc22241, nc22242, nc22243, 
        nc22244, nc22245, nc22246, nc22247, \R_DATA_TEMPR17[35] , 
        \R_DATA_TEMPR17[34] }), .B_DOUT({nc22248, nc22249, nc22250, 
        nc22251, nc22252, nc22253, nc22254, nc22255, nc22256, nc22257, 
        nc22258, nc22259, nc22260, nc22261, nc22262, nc22263, nc22264, 
        nc22265, nc22266, nc22267}), .DB_DETECT(\DB_DETECT[17][17] ), 
        .SB_CORRECT(\SB_CORRECT[17][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_137 (.A(\R_DATA_TEMPR16[33] ), .B(\R_DATA_TEMPR17[33] ), 
        .C(\R_DATA_TEMPR18[33] ), .D(\R_DATA_TEMPR19[33] ), .Y(
        OR4_137_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C16 (.A_DOUT({
        nc22268, nc22269, nc22270, nc22271, nc22272, nc22273, nc22274, 
        nc22275, nc22276, nc22277, nc22278, nc22279, nc22280, nc22281, 
        nc22282, nc22283, nc22284, nc22285, \R_DATA_TEMPR6[33] , 
        \R_DATA_TEMPR6[32] }), .B_DOUT({nc22286, nc22287, nc22288, 
        nc22289, nc22290, nc22291, nc22292, nc22293, nc22294, nc22295, 
        nc22296, nc22297, nc22298, nc22299, nc22300, nc22301, nc22302, 
        nc22303, nc22304, nc22305}), .DB_DETECT(\DB_DETECT[6][16] ), 
        .SB_CORRECT(\SB_CORRECT[6][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C11 (.A_DOUT({
        nc22306, nc22307, nc22308, nc22309, nc22310, nc22311, nc22312, 
        nc22313, nc22314, nc22315, nc22316, nc22317, nc22318, nc22319, 
        nc22320, nc22321, nc22322, nc22323, \R_DATA_TEMPR3[23] , 
        \R_DATA_TEMPR3[22] }), .B_DOUT({nc22324, nc22325, nc22326, 
        nc22327, nc22328, nc22329, nc22330, nc22331, nc22332, nc22333, 
        nc22334, nc22335, nc22336, nc22337, nc22338, nc22339, nc22340, 
        nc22341, nc22342, nc22343}), .DB_DETECT(\DB_DETECT[3][11] ), 
        .SB_CORRECT(\SB_CORRECT[3][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_342 (.A(OR4_286_Y), .B(OR4_359_Y), .C(OR4_30_Y), .D(
        OR4_300_Y), .Y(OR4_342_Y));
    OR4 OR4_359 (.A(\R_DATA_TEMPR4[14] ), .B(\R_DATA_TEMPR5[14] ), .C(
        \R_DATA_TEMPR6[14] ), .D(\R_DATA_TEMPR7[14] ), .Y(OR4_359_Y));
    OR4 OR4_14 (.A(OR4_354_Y), .B(OR4_272_Y), .C(OR4_358_Y), .D(
        OR4_148_Y), .Y(OR4_14_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C19 (.A_DOUT({
        nc22344, nc22345, nc22346, nc22347, nc22348, nc22349, nc22350, 
        nc22351, nc22352, nc22353, nc22354, nc22355, nc22356, nc22357, 
        nc22358, nc22359, nc22360, nc22361, \R_DATA_TEMPR5[39] , 
        \R_DATA_TEMPR5[38] }), .B_DOUT({nc22362, nc22363, nc22364, 
        nc22365, nc22366, nc22367, nc22368, nc22369, nc22370, nc22371, 
        nc22372, nc22373, nc22374, nc22375, nc22376, nc22377, nc22378, 
        nc22379, nc22380, nc22381}), .DB_DETECT(\DB_DETECT[5][19] ), 
        .SB_CORRECT(\SB_CORRECT[5][19] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][19] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[39], W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[19]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C6 (.A_DOUT({nc22382, 
        nc22383, nc22384, nc22385, nc22386, nc22387, nc22388, nc22389, 
        nc22390, nc22391, nc22392, nc22393, nc22394, nc22395, nc22396, 
        nc22397, nc22398, nc22399, \R_DATA_TEMPR6[13] , 
        \R_DATA_TEMPR6[12] }), .B_DOUT({nc22400, nc22401, nc22402, 
        nc22403, nc22404, nc22405, nc22406, nc22407, nc22408, nc22409, 
        nc22410, nc22411, nc22412, nc22413, nc22414, nc22415, nc22416, 
        nc22417, nc22418, nc22419}), .DB_DETECT(\DB_DETECT[6][6] ), 
        .SB_CORRECT(\SB_CORRECT[6][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[6][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C12 (.A_DOUT({
        nc22420, nc22421, nc22422, nc22423, nc22424, nc22425, nc22426, 
        nc22427, nc22428, nc22429, nc22430, nc22431, nc22432, nc22433, 
        nc22434, nc22435, nc22436, nc22437, \R_DATA_TEMPR16[25] , 
        \R_DATA_TEMPR16[24] }), .B_DOUT({nc22438, nc22439, nc22440, 
        nc22441, nc22442, nc22443, nc22444, nc22445, nc22446, nc22447, 
        nc22448, nc22449, nc22450, nc22451, nc22452, nc22453, nc22454, 
        nc22455, nc22456, nc22457}), .DB_DETECT(\DB_DETECT[16][12] ), 
        .SB_CORRECT(\SB_CORRECT[16][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[16][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C11 (.A_DOUT({
        nc22458, nc22459, nc22460, nc22461, nc22462, nc22463, nc22464, 
        nc22465, nc22466, nc22467, nc22468, nc22469, nc22470, nc22471, 
        nc22472, nc22473, nc22474, nc22475, \R_DATA_TEMPR26[23] , 
        \R_DATA_TEMPR26[22] }), .B_DOUT({nc22476, nc22477, nc22478, 
        nc22479, nc22480, nc22481, nc22482, nc22483, nc22484, nc22485, 
        nc22486, nc22487, nc22488, nc22489, nc22490, nc22491, nc22492, 
        nc22493, nc22494, nc22495}), .DB_DETECT(\DB_DETECT[26][11] ), 
        .SB_CORRECT(\SB_CORRECT[26][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_18 (.A(\R_DATA_TEMPR20[38] ), .B(\R_DATA_TEMPR21[38] ), .Y(
        OR2_18_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C2 (.A_DOUT({
        nc22496, nc22497, nc22498, nc22499, nc22500, nc22501, nc22502, 
        nc22503, nc22504, nc22505, nc22506, nc22507, nc22508, nc22509, 
        nc22510, nc22511, nc22512, nc22513, \R_DATA_TEMPR26[5] , 
        \R_DATA_TEMPR26[4] }), .B_DOUT({nc22514, nc22515, nc22516, 
        nc22517, nc22518, nc22519, nc22520, nc22521, nc22522, nc22523, 
        nc22524, nc22525, nc22526, nc22527, nc22528, nc22529, nc22530, 
        nc22531, nc22532, nc22533}), .DB_DETECT(\DB_DETECT[26][2] ), 
        .SB_CORRECT(\SB_CORRECT[26][2] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][2] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[5], W_DATA[4]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C7 (.A_DOUT({
        nc22534, nc22535, nc22536, nc22537, nc22538, nc22539, nc22540, 
        nc22541, nc22542, nc22543, nc22544, nc22545, nc22546, nc22547, 
        nc22548, nc22549, nc22550, nc22551, \R_DATA_TEMPR26[15] , 
        \R_DATA_TEMPR26[14] }), .B_DOUT({nc22552, nc22553, nc22554, 
        nc22555, nc22556, nc22557, nc22558, nc22559, nc22560, nc22561, 
        nc22562, nc22563, nc22564, nc22565, nc22566, nc22567, nc22568, 
        nc22569, nc22570, nc22571}), .DB_DETECT(\DB_DETECT[26][7] ), 
        .SB_CORRECT(\SB_CORRECT[26][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[26][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_291 (.A(\R_DATA_TEMPR12[29] ), .B(\R_DATA_TEMPR13[29] ), 
        .C(\R_DATA_TEMPR14[29] ), .D(\R_DATA_TEMPR15[29] ), .Y(
        OR4_291_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C3 (.A_DOUT({nc22572, 
        nc22573, nc22574, nc22575, nc22576, nc22577, nc22578, nc22579, 
        nc22580, nc22581, nc22582, nc22583, nc22584, nc22585, nc22586, 
        nc22587, nc22588, nc22589, \R_DATA_TEMPR3[7] , 
        \R_DATA_TEMPR3[6] }), .B_DOUT({nc22590, nc22591, nc22592, 
        nc22593, nc22594, nc22595, nc22596, nc22597, nc22598, nc22599, 
        nc22600, nc22601, nc22602, nc22603, nc22604, nc22605, nc22606, 
        nc22607, nc22608, nc22609}), .DB_DETECT(\DB_DETECT[3][3] ), 
        .SB_CORRECT(\SB_CORRECT[3][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[3][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C14 (.A_DOUT({
        nc22610, nc22611, nc22612, nc22613, nc22614, nc22615, nc22616, 
        nc22617, nc22618, nc22619, nc22620, nc22621, nc22622, nc22623, 
        nc22624, nc22625, nc22626, nc22627, \R_DATA_TEMPR23[29] , 
        \R_DATA_TEMPR23[28] }), .B_DOUT({nc22628, nc22629, nc22630, 
        nc22631, nc22632, nc22633, nc22634, nc22635, nc22636, nc22637, 
        nc22638, nc22639, nc22640, nc22641, nc22642, nc22643, nc22644, 
        nc22645, nc22646, nc22647}), .DB_DETECT(\DB_DETECT[23][14] ), 
        .SB_CORRECT(\SB_CORRECT[23][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C12 (.A_DOUT({
        nc22648, nc22649, nc22650, nc22651, nc22652, nc22653, nc22654, 
        nc22655, nc22656, nc22657, nc22658, nc22659, nc22660, nc22661, 
        nc22662, nc22663, nc22664, nc22665, \R_DATA_TEMPR24[25] , 
        \R_DATA_TEMPR24[24] }), .B_DOUT({nc22666, nc22667, nc22668, 
        nc22669, nc22670, nc22671, nc22672, nc22673, nc22674, nc22675, 
        nc22676, nc22677, nc22678, nc22679, nc22680, nc22681, nc22682, 
        nc22683, nc22684, nc22685}), .DB_DETECT(\DB_DETECT[24][12] ), 
        .SB_CORRECT(\SB_CORRECT[24][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_234 (.A(\R_DATA_TEMPR8[2] ), .B(\R_DATA_TEMPR9[2] ), .C(
        \R_DATA_TEMPR10[2] ), .D(\R_DATA_TEMPR11[2] ), .Y(OR4_234_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C10 (.A_DOUT({
        nc22686, nc22687, nc22688, nc22689, nc22690, nc22691, nc22692, 
        nc22693, nc22694, nc22695, nc22696, nc22697, nc22698, nc22699, 
        nc22700, nc22701, nc22702, nc22703, \R_DATA_TEMPR24[21] , 
        \R_DATA_TEMPR24[20] }), .B_DOUT({nc22704, nc22705, nc22706, 
        nc22707, nc22708, nc22709, nc22710, nc22711, nc22712, nc22713, 
        nc22714, nc22715, nc22716, nc22717, nc22718, nc22719, nc22720, 
        nc22721, nc22722, nc22723}), .DB_DETECT(\DB_DETECT[24][10] ), 
        .SB_CORRECT(\SB_CORRECT[24][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C13 (.A_DOUT({
        nc22724, nc22725, nc22726, nc22727, nc22728, nc22729, nc22730, 
        nc22731, nc22732, nc22733, nc22734, nc22735, nc22736, nc22737, 
        nc22738, nc22739, nc22740, nc22741, \R_DATA_TEMPR31[27] , 
        \R_DATA_TEMPR31[26] }), .B_DOUT({nc22742, nc22743, nc22744, 
        nc22745, nc22746, nc22747, nc22748, nc22749, nc22750, nc22751, 
        nc22752, nc22753, nc22754, nc22755, nc22756, nc22757, nc22758, 
        nc22759, nc22760, nc22761}), .DB_DETECT(\DB_DETECT[31][13] ), 
        .SB_CORRECT(\SB_CORRECT[31][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C15 (.A_DOUT({
        nc22762, nc22763, nc22764, nc22765, nc22766, nc22767, nc22768, 
        nc22769, nc22770, nc22771, nc22772, nc22773, nc22774, nc22775, 
        nc22776, nc22777, nc22778, nc22779, \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR4[30] }), .B_DOUT({nc22780, nc22781, nc22782, 
        nc22783, nc22784, nc22785, nc22786, nc22787, nc22788, nc22789, 
        nc22790, nc22791, nc22792, nc22793, nc22794, nc22795, nc22796, 
        nc22797, nc22798, nc22799}), .DB_DETECT(\DB_DETECT[4][15] ), 
        .SB_CORRECT(\SB_CORRECT[4][15] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][15] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[31], W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[15]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C6 (.A_DOUT({
        nc22800, nc22801, nc22802, nc22803, nc22804, nc22805, nc22806, 
        nc22807, nc22808, nc22809, nc22810, nc22811, nc22812, nc22813, 
        nc22814, nc22815, nc22816, nc22817, \R_DATA_TEMPR12[13] , 
        \R_DATA_TEMPR12[12] }), .B_DOUT({nc22818, nc22819, nc22820, 
        nc22821, nc22822, nc22823, nc22824, nc22825, nc22826, nc22827, 
        nc22828, nc22829, nc22830, nc22831, nc22832, nc22833, nc22834, 
        nc22835, nc22836, nc22837}), .DB_DETECT(\DB_DETECT[12][6] ), 
        .SB_CORRECT(\SB_CORRECT[12][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_90 (.A(\R_DATA_TEMPR8[6] ), .B(\R_DATA_TEMPR9[6] ), .C(
        \R_DATA_TEMPR10[6] ), .D(\R_DATA_TEMPR11[6] ), .Y(OR4_90_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C7 (.A_DOUT({
        nc22838, nc22839, nc22840, nc22841, nc22842, nc22843, nc22844, 
        nc22845, nc22846, nc22847, nc22848, nc22849, nc22850, nc22851, 
        nc22852, nc22853, nc22854, nc22855, \R_DATA_TEMPR22[15] , 
        \R_DATA_TEMPR22[14] }), .B_DOUT({nc22856, nc22857, nc22858, 
        nc22859, nc22860, nc22861, nc22862, nc22863, nc22864, nc22865, 
        nc22866, nc22867, nc22868, nc22869, nc22870, nc22871, nc22872, 
        nc22873, nc22874, nc22875}), .DB_DETECT(\DB_DETECT[22][7] ), 
        .SB_CORRECT(\SB_CORRECT[22][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[22][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C12 (.A_DOUT({
        nc22876, nc22877, nc22878, nc22879, nc22880, nc22881, nc22882, 
        nc22883, nc22884, nc22885, nc22886, nc22887, nc22888, nc22889, 
        nc22890, nc22891, nc22892, nc22893, \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR1[24] }), .B_DOUT({nc22894, nc22895, nc22896, 
        nc22897, nc22898, nc22899, nc22900, nc22901, nc22902, nc22903, 
        nc22904, nc22905, nc22906, nc22907, nc22908, nc22909, nc22910, 
        nc22911, nc22912, nc22913}), .DB_DETECT(\DB_DETECT[1][12] ), 
        .SB_CORRECT(\SB_CORRECT[1][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[1][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C8 (.A_DOUT({nc22914, 
        nc22915, nc22916, nc22917, nc22918, nc22919, nc22920, nc22921, 
        nc22922, nc22923, nc22924, nc22925, nc22926, nc22927, nc22928, 
        nc22929, nc22930, nc22931, \R_DATA_TEMPR8[17] , 
        \R_DATA_TEMPR8[16] }), .B_DOUT({nc22932, nc22933, nc22934, 
        nc22935, nc22936, nc22937, nc22938, nc22939, nc22940, nc22941, 
        nc22942, nc22943, nc22944, nc22945, nc22946, nc22947, nc22948, 
        nc22949, nc22950, nc22951}), .DB_DETECT(\DB_DETECT[8][8] ), 
        .SB_CORRECT(\SB_CORRECT[8][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C12 (.A_DOUT({
        nc22952, nc22953, nc22954, nc22955, nc22956, nc22957, nc22958, 
        nc22959, nc22960, nc22961, nc22962, nc22963, nc22964, nc22965, 
        nc22966, nc22967, nc22968, nc22969, \R_DATA_TEMPR25[25] , 
        \R_DATA_TEMPR25[24] }), .B_DOUT({nc22970, nc22971, nc22972, 
        nc22973, nc22974, nc22975, nc22976, nc22977, nc22978, nc22979, 
        nc22980, nc22981, nc22982, nc22983, nc22984, nc22985, nc22986, 
        nc22987, nc22988, nc22989}), .DB_DETECT(\DB_DETECT[25][12] ), 
        .SB_CORRECT(\SB_CORRECT[25][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_46 (.A(\R_DATA_TEMPR16[0] ), .B(\R_DATA_TEMPR17[0] ), .C(
        \R_DATA_TEMPR18[0] ), .D(\R_DATA_TEMPR19[0] ), .Y(OR4_46_Y));
    OR4 OR4_97 (.A(OR4_313_Y), .B(OR2_22_Y), .C(\R_DATA_TEMPR22[25] ), 
        .D(\R_DATA_TEMPR23[25] ), .Y(OR4_97_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C10 (.A_DOUT({
        nc22990, nc22991, nc22992, nc22993, nc22994, nc22995, nc22996, 
        nc22997, nc22998, nc22999, nc23000, nc23001, nc23002, nc23003, 
        nc23004, nc23005, nc23006, nc23007, \R_DATA_TEMPR25[21] , 
        \R_DATA_TEMPR25[20] }), .B_DOUT({nc23008, nc23009, nc23010, 
        nc23011, nc23012, nc23013, nc23014, nc23015, nc23016, nc23017, 
        nc23018, nc23019, nc23020, nc23021, nc23022, nc23023, nc23024, 
        nc23025, nc23026, nc23027}), .DB_DETECT(\DB_DETECT[25][10] ), 
        .SB_CORRECT(\SB_CORRECT[25][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C5 (.A_DOUT({nc23028, 
        nc23029, nc23030, nc23031, nc23032, nc23033, nc23034, nc23035, 
        nc23036, nc23037, nc23038, nc23039, nc23040, nc23041, nc23042, 
        nc23043, nc23044, nc23045, \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR8[10] }), .B_DOUT({nc23046, nc23047, nc23048, 
        nc23049, nc23050, nc23051, nc23052, nc23053, nc23054, nc23055, 
        nc23056, nc23057, nc23058, nc23059, nc23060, nc23061, nc23062, 
        nc23063, nc23064, nc23065}), .DB_DETECT(\DB_DETECT[8][5] ), 
        .SB_CORRECT(\SB_CORRECT[8][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[6]  (.A(OR4_82_Y), .B(OR4_251_Y), .C(OR4_11_Y), .D(
        OR4_55_Y), .Y(R_DATA[6]));
    OR4 OR4_63 (.A(\R_DATA_TEMPR24[16] ), .B(\R_DATA_TEMPR25[16] ), .C(
        \R_DATA_TEMPR26[16] ), .D(\R_DATA_TEMPR27[16] ), .Y(OR4_63_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C13 (.A_DOUT({
        nc23066, nc23067, nc23068, nc23069, nc23070, nc23071, nc23072, 
        nc23073, nc23074, nc23075, nc23076, nc23077, nc23078, nc23079, 
        nc23080, nc23081, nc23082, nc23083, \R_DATA_TEMPR10[27] , 
        \R_DATA_TEMPR10[26] }), .B_DOUT({nc23084, nc23085, nc23086, 
        nc23087, nc23088, nc23089, nc23090, nc23091, nc23092, nc23093, 
        nc23094, nc23095, nc23096, nc23097, nc23098, nc23099, nc23100, 
        nc23101, nc23102, nc23103}), .DB_DETECT(\DB_DETECT[10][13] ), 
        .SB_CORRECT(\SB_CORRECT[10][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[10][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_217 (.A(\R_DATA_TEMPR8[26] ), .B(\R_DATA_TEMPR9[26] ), .C(
        \R_DATA_TEMPR10[26] ), .D(\R_DATA_TEMPR11[26] ), .Y(OR4_217_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C16 (.A_DOUT({
        nc23104, nc23105, nc23106, nc23107, nc23108, nc23109, nc23110, 
        nc23111, nc23112, nc23113, nc23114, nc23115, nc23116, nc23117, 
        nc23118, nc23119, nc23120, nc23121, \R_DATA_TEMPR14[33] , 
        \R_DATA_TEMPR14[32] }), .B_DOUT({nc23122, nc23123, nc23124, 
        nc23125, nc23126, nc23127, nc23128, nc23129, nc23130, nc23131, 
        nc23132, nc23133, nc23134, nc23135, nc23136, nc23137, nc23138, 
        nc23139, nc23140, nc23141}), .DB_DETECT(\DB_DETECT[14][16] ), 
        .SB_CORRECT(\SB_CORRECT[14][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_304 (.A(\R_DATA_TEMPR28[19] ), .B(\R_DATA_TEMPR29[19] ), 
        .C(\R_DATA_TEMPR30[19] ), .D(\R_DATA_TEMPR31[19] ), .Y(
        OR4_304_Y));
    OR4 OR4_240 (.A(\R_DATA_TEMPR16[2] ), .B(\R_DATA_TEMPR17[2] ), .C(
        \R_DATA_TEMPR18[2] ), .D(\R_DATA_TEMPR19[2] ), .Y(OR4_240_Y));
    OR4 OR4_117 (.A(OR4_254_Y), .B(OR4_16_Y), .C(OR4_166_Y), .D(
        OR4_322_Y), .Y(OR4_117_Y));
    OR4 OR4_335 (.A(\R_DATA_TEMPR12[37] ), .B(\R_DATA_TEMPR13[37] ), 
        .C(\R_DATA_TEMPR14[37] ), .D(\R_DATA_TEMPR15[37] ), .Y(
        OR4_335_Y));
    OR4 \OR4_R_DATA[1]  (.A(OR4_292_Y), .B(OR4_334_Y), .C(OR4_236_Y), 
        .D(OR4_188_Y), .Y(R_DATA[1]));
    OR4 OR4_101 (.A(\R_DATA_TEMPR16[7] ), .B(\R_DATA_TEMPR17[7] ), .C(
        \R_DATA_TEMPR18[7] ), .D(\R_DATA_TEMPR19[7] ), .Y(OR4_101_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C16 (.A_DOUT({
        nc23142, nc23143, nc23144, nc23145, nc23146, nc23147, nc23148, 
        nc23149, nc23150, nc23151, nc23152, nc23153, nc23154, nc23155, 
        nc23156, nc23157, nc23158, nc23159, \R_DATA_TEMPR15[33] , 
        \R_DATA_TEMPR15[32] }), .B_DOUT({nc23160, nc23161, nc23162, 
        nc23163, nc23164, nc23165, nc23166, nc23167, nc23168, nc23169, 
        nc23170, nc23171, nc23172, nc23173, nc23174, nc23175, nc23176, 
        nc23177, nc23178, nc23179}), .DB_DETECT(\DB_DETECT[15][16] ), 
        .SB_CORRECT(\SB_CORRECT[15][16] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][16] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[33], W_DATA[32]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[16]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C5 (.A_DOUT({
        nc23180, nc23181, nc23182, nc23183, nc23184, nc23185, nc23186, 
        nc23187, nc23188, nc23189, nc23190, nc23191, nc23192, nc23193, 
        nc23194, nc23195, nc23196, nc23197, \R_DATA_TEMPR31[11] , 
        \R_DATA_TEMPR31[10] }), .B_DOUT({nc23198, nc23199, nc23200, 
        nc23201, nc23202, nc23203, nc23204, nc23205, nc23206, nc23207, 
        nc23208, nc23209, nc23210, nc23211, nc23212, nc23213, nc23214, 
        nc23215, nc23216, nc23217}), .DB_DETECT(\DB_DETECT[31][5] ), 
        .SB_CORRECT(\SB_CORRECT[31][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C11 (.A_DOUT({
        nc23218, nc23219, nc23220, nc23221, nc23222, nc23223, nc23224, 
        nc23225, nc23226, nc23227, nc23228, nc23229, nc23230, nc23231, 
        nc23232, nc23233, nc23234, nc23235, \R_DATA_TEMPR11[23] , 
        \R_DATA_TEMPR11[22] }), .B_DOUT({nc23236, nc23237, nc23238, 
        nc23239, nc23240, nc23241, nc23242, nc23243, nc23244, nc23245, 
        nc23246, nc23247, nc23248, nc23249, nc23250, nc23251, nc23252, 
        nc23253, nc23254, nc23255}), .DB_DETECT(\DB_DETECT[11][11] ), 
        .SB_CORRECT(\SB_CORRECT[11][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[11][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C17 (.A_DOUT({
        nc23256, nc23257, nc23258, nc23259, nc23260, nc23261, nc23262, 
        nc23263, nc23264, nc23265, nc23266, nc23267, nc23268, nc23269, 
        nc23270, nc23271, nc23272, nc23273, \R_DATA_TEMPR12[35] , 
        \R_DATA_TEMPR12[34] }), .B_DOUT({nc23274, nc23275, nc23276, 
        nc23277, nc23278, nc23279, nc23280, nc23281, nc23282, nc23283, 
        nc23284, nc23285, nc23286, nc23287, nc23288, nc23289, nc23290, 
        nc23291, nc23292, nc23293}), .DB_DETECT(\DB_DETECT[12][17] ), 
        .SB_CORRECT(\SB_CORRECT[12][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[12][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_171 (.A(\R_DATA_TEMPR24[10] ), .B(\R_DATA_TEMPR25[10] ), 
        .C(\R_DATA_TEMPR26[10] ), .D(\R_DATA_TEMPR27[10] ), .Y(
        OR4_171_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C3 (.A_DOUT({
        nc23294, nc23295, nc23296, nc23297, nc23298, nc23299, nc23300, 
        nc23301, nc23302, nc23303, nc23304, nc23305, nc23306, nc23307, 
        nc23308, nc23309, nc23310, nc23311, \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR24[6] }), .B_DOUT({nc23312, nc23313, nc23314, 
        nc23315, nc23316, nc23317, nc23318, nc23319, nc23320, nc23321, 
        nc23322, nc23323, nc23324, nc23325, nc23326, nc23327, nc23328, 
        nc23329, nc23330, nc23331}), .DB_DETECT(\DB_DETECT[24][3] ), 
        .SB_CORRECT(\SB_CORRECT[24][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C17 (.A_DOUT({
        nc23332, nc23333, nc23334, nc23335, nc23336, nc23337, nc23338, 
        nc23339, nc23340, nc23341, nc23342, nc23343, nc23344, nc23345, 
        nc23346, nc23347, nc23348, nc23349, \R_DATA_TEMPR20[35] , 
        \R_DATA_TEMPR20[34] }), .B_DOUT({nc23350, nc23351, nc23352, 
        nc23353, nc23354, nc23355, nc23356, nc23357, nc23358, nc23359, 
        nc23360, nc23361, nc23362, nc23363, nc23364, nc23365, nc23366, 
        nc23367, nc23368, nc23369}), .DB_DETECT(\DB_DETECT[20][17] ), 
        .SB_CORRECT(\SB_CORRECT[20][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C9 (.A_DOUT({
        nc23370, nc23371, nc23372, nc23373, nc23374, nc23375, nc23376, 
        nc23377, nc23378, nc23379, nc23380, nc23381, nc23382, nc23383, 
        nc23384, nc23385, nc23386, nc23387, \R_DATA_TEMPR20[19] , 
        \R_DATA_TEMPR20[18] }), .B_DOUT({nc23388, nc23389, nc23390, 
        nc23391, nc23392, nc23393, nc23394, nc23395, nc23396, nc23397, 
        nc23398, nc23399, nc23400, nc23401, nc23402, nc23403, nc23404, 
        nc23405, nc23406, nc23407}), .DB_DETECT(\DB_DETECT[20][9] ), 
        .SB_CORRECT(\SB_CORRECT[20][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_214 (.A(OR4_235_Y), .B(OR2_21_Y), .C(\R_DATA_TEMPR22[8] ), 
        .D(\R_DATA_TEMPR23[8] ), .Y(OR4_214_Y));
    OR4 OR4_246 (.A(OR4_57_Y), .B(OR4_317_Y), .C(OR4_333_Y), .D(
        OR4_31_Y), .Y(OR4_246_Y));
    OR4 OR4_221 (.A(\R_DATA_TEMPR4[3] ), .B(\R_DATA_TEMPR5[3] ), .C(
        \R_DATA_TEMPR6[3] ), .D(\R_DATA_TEMPR7[3] ), .Y(OR4_221_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C9 (.A_DOUT({nc23408, 
        nc23409, nc23410, nc23411, nc23412, nc23413, nc23414, nc23415, 
        nc23416, nc23417, nc23418, nc23419, nc23420, nc23421, nc23422, 
        nc23423, nc23424, nc23425, \R_DATA_TEMPR0[19] , 
        \R_DATA_TEMPR0[18] }), .B_DOUT({nc23426, nc23427, nc23428, 
        nc23429, nc23430, nc23431, nc23432, nc23433, nc23434, nc23435, 
        nc23436, nc23437, nc23438, nc23439, nc23440, nc23441, nc23442, 
        nc23443, nc23444, nc23445}), .DB_DETECT(\DB_DETECT[0][9] ), 
        .SB_CORRECT(\SB_CORRECT[0][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_74 (.A(\R_DATA_TEMPR16[28] ), .B(\R_DATA_TEMPR17[28] ), .C(
        \R_DATA_TEMPR18[28] ), .D(\R_DATA_TEMPR19[28] ), .Y(OR4_74_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[6]  (.A(CFG2_7_Y), .B(
        W_ADDR[17]), .C(W_EN), .Y(\BLKX2[6] ));
    OR4 OR4_61 (.A(OR4_165_Y), .B(OR2_19_Y), .C(\R_DATA_TEMPR22[31] ), 
        .D(\R_DATA_TEMPR23[31] ), .Y(OR4_61_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C6 (.A_DOUT({
        nc23446, nc23447, nc23448, nc23449, nc23450, nc23451, nc23452, 
        nc23453, nc23454, nc23455, nc23456, nc23457, nc23458, nc23459, 
        nc23460, nc23461, nc23462, nc23463, \R_DATA_TEMPR20[13] , 
        \R_DATA_TEMPR20[12] }), .B_DOUT({nc23464, nc23465, nc23466, 
        nc23467, nc23468, nc23469, nc23470, nc23471, nc23472, nc23473, 
        nc23474, nc23475, nc23476, nc23477, nc23478, nc23479, nc23480, 
        nc23481, nc23482, nc23483}), .DB_DETECT(\DB_DETECT[20][6] ), 
        .SB_CORRECT(\SB_CORRECT[20][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C12 (.A_DOUT({
        nc23484, nc23485, nc23486, nc23487, nc23488, nc23489, nc23490, 
        nc23491, nc23492, nc23493, nc23494, nc23495, nc23496, nc23497, 
        nc23498, nc23499, nc23500, nc23501, \R_DATA_TEMPR8[25] , 
        \R_DATA_TEMPR8[24] }), .B_DOUT({nc23502, nc23503, nc23504, 
        nc23505, nc23506, nc23507, nc23508, nc23509, nc23510, nc23511, 
        nc23512, nc23513, nc23514, nc23515, nc23516, nc23517, nc23518, 
        nc23519, nc23520, nc23521}), .DB_DETECT(\DB_DETECT[8][12] ), 
        .SB_CORRECT(\SB_CORRECT[8][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[8][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C5 (.A_DOUT({nc23522, 
        nc23523, nc23524, nc23525, nc23526, nc23527, nc23528, nc23529, 
        nc23530, nc23531, nc23532, nc23533, nc23534, nc23535, nc23536, 
        nc23537, nc23538, nc23539, \R_DATA_TEMPR7[11] , 
        \R_DATA_TEMPR7[10] }), .B_DOUT({nc23540, nc23541, nc23542, 
        nc23543, nc23544, nc23545, nc23546, nc23547, nc23548, nc23549, 
        nc23550, nc23551, nc23552, nc23553, nc23554, nc23555, nc23556, 
        nc23557, nc23558, nc23559}), .DB_DETECT(\DB_DETECT[7][5] ), 
        .SB_CORRECT(\SB_CORRECT[7][5] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][5] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[11], W_DATA[10]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[5]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C13 (.A_DOUT({
        nc23560, nc23561, nc23562, nc23563, nc23564, nc23565, nc23566, 
        nc23567, nc23568, nc23569, nc23570, nc23571, nc23572, nc23573, 
        nc23574, nc23575, nc23576, nc23577, \R_DATA_TEMPR9[27] , 
        \R_DATA_TEMPR9[26] }), .B_DOUT({nc23578, nc23579, nc23580, 
        nc23581, nc23582, nc23583, nc23584, nc23585, nc23586, nc23587, 
        nc23588, nc23589, nc23590, nc23591, nc23592, nc23593, nc23594, 
        nc23595, nc23596, nc23597}), .DB_DETECT(\DB_DETECT[9][13] ), 
        .SB_CORRECT(\SB_CORRECT[9][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[9][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_315 (.A(\R_DATA_TEMPR4[9] ), .B(\R_DATA_TEMPR5[9] ), .C(
        \R_DATA_TEMPR6[9] ), .D(\R_DATA_TEMPR7[9] ), .Y(OR4_315_Y));
    OR2 OR2_5 (.A(\R_DATA_TEMPR20[5] ), .B(\R_DATA_TEMPR21[5] ), .Y(
        OR2_5_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C13 (.A_DOUT({
        nc23598, nc23599, nc23600, nc23601, nc23602, nc23603, nc23604, 
        nc23605, nc23606, nc23607, nc23608, nc23609, nc23610, nc23611, 
        nc23612, nc23613, nc23614, nc23615, \R_DATA_TEMPR14[27] , 
        \R_DATA_TEMPR14[26] }), .B_DOUT({nc23616, nc23617, nc23618, 
        nc23619, nc23620, nc23621, nc23622, nc23623, nc23624, nc23625, 
        nc23626, nc23627, nc23628, nc23629, nc23630, nc23631, nc23632, 
        nc23633, nc23634, nc23635}), .DB_DETECT(\DB_DETECT[14][13] ), 
        .SB_CORRECT(\SB_CORRECT[14][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_40 (.A(OR4_76_Y), .B(OR4_276_Y), .C(OR4_45_Y), .D(
        OR4_219_Y), .Y(OR4_40_Y));
    OR4 OR4_166 (.A(\R_DATA_TEMPR8[19] ), .B(\R_DATA_TEMPR9[19] ), .C(
        \R_DATA_TEMPR10[19] ), .D(\R_DATA_TEMPR11[19] ), .Y(OR4_166_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C6 (.A_DOUT({nc23636, 
        nc23637, nc23638, nc23639, nc23640, nc23641, nc23642, nc23643, 
        nc23644, nc23645, nc23646, nc23647, nc23648, nc23649, nc23650, 
        nc23651, nc23652, nc23653, \R_DATA_TEMPR5[13] , 
        \R_DATA_TEMPR5[12] }), .B_DOUT({nc23654, nc23655, nc23656, 
        nc23657, nc23658, nc23659, nc23660, nc23661, nc23662, nc23663, 
        nc23664, nc23665, nc23666, nc23667, nc23668, nc23669, nc23670, 
        nc23671, nc23672, nc23673}), .DB_DETECT(\DB_DETECT[5][6] ), 
        .SB_CORRECT(\SB_CORRECT[5][6] ), .ACCESS_BUSY(
        \ACCESS_BUSY[5][6] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[13], W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C13 (.A_DOUT({
        nc23674, nc23675, nc23676, nc23677, nc23678, nc23679, nc23680, 
        nc23681, nc23682, nc23683, nc23684, nc23685, nc23686, nc23687, 
        nc23688, nc23689, nc23690, nc23691, \R_DATA_TEMPR23[27] , 
        \R_DATA_TEMPR23[26] }), .B_DOUT({nc23692, nc23693, nc23694, 
        nc23695, nc23696, nc23697, nc23698, nc23699, nc23700, nc23701, 
        nc23702, nc23703, nc23704, nc23705, nc23706, nc23707, nc23708, 
        nc23709, nc23710, nc23711}), .DB_DETECT(\DB_DETECT[23][13] ), 
        .SB_CORRECT(\SB_CORRECT[23][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[23][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C14 (.A_DOUT({
        nc23712, nc23713, nc23714, nc23715, nc23716, nc23717, nc23718, 
        nc23719, nc23720, nc23721, nc23722, nc23723, nc23724, nc23725, 
        nc23726, nc23727, nc23728, nc23729, \R_DATA_TEMPR20[29] , 
        \R_DATA_TEMPR20[28] }), .B_DOUT({nc23730, nc23731, nc23732, 
        nc23733, nc23734, nc23735, nc23736, nc23737, nc23738, nc23739, 
        nc23740, nc23741, nc23742, nc23743, nc23744, nc23745, nc23746, 
        nc23747, nc23748, nc23749}), .DB_DETECT(\DB_DETECT[20][14] ), 
        .SB_CORRECT(\SB_CORRECT[20][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[20][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_47 (.A(\R_DATA_TEMPR0[8] ), .B(\R_DATA_TEMPR1[8] ), .C(
        \R_DATA_TEMPR2[8] ), .D(\R_DATA_TEMPR3[8] ), .Y(OR4_47_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C14 (.A_DOUT({
        nc23750, nc23751, nc23752, nc23753, nc23754, nc23755, nc23756, 
        nc23757, nc23758, nc23759, nc23760, nc23761, nc23762, nc23763, 
        nc23764, nc23765, nc23766, nc23767, \R_DATA_TEMPR18[29] , 
        \R_DATA_TEMPR18[28] }), .B_DOUT({nc23768, nc23769, nc23770, 
        nc23771, nc23772, nc23773, nc23774, nc23775, nc23776, nc23777, 
        nc23778, nc23779, nc23780, nc23781, nc23782, nc23783, nc23784, 
        nc23785, nc23786, nc23787}), .DB_DETECT(\DB_DETECT[18][14] ), 
        .SB_CORRECT(\SB_CORRECT[18][14] ), .ACCESS_BUSY(
        \ACCESS_BUSY[18][14] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[29], W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[14]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0 (.A_DOUT({nc23788, 
        nc23789, nc23790, nc23791, nc23792, nc23793, nc23794, nc23795, 
        nc23796, nc23797, nc23798, nc23799, nc23800, nc23801, nc23802, 
        nc23803, nc23804, nc23805, \R_DATA_TEMPR7[1] , 
        \R_DATA_TEMPR7[0] }), .B_DOUT({nc23806, nc23807, nc23808, 
        nc23809, nc23810, nc23811, nc23812, nc23813, nc23814, nc23815, 
        nc23816, nc23817, nc23818, nc23819, nc23820, nc23821, nc23822, 
        nc23823, nc23824, nc23825}), .DB_DETECT(\DB_DETECT[7][0] ), 
        .SB_CORRECT(\SB_CORRECT[7][0] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][0] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C13 (.A_DOUT({
        nc23826, nc23827, nc23828, nc23829, nc23830, nc23831, nc23832, 
        nc23833, nc23834, nc23835, nc23836, nc23837, nc23838, nc23839, 
        nc23840, nc23841, nc23842, nc23843, \R_DATA_TEMPR15[27] , 
        \R_DATA_TEMPR15[26] }), .B_DOUT({nc23844, nc23845, nc23846, 
        nc23847, nc23848, nc23849, nc23850, nc23851, nc23852, nc23853, 
        nc23854, nc23855, nc23856, nc23857, nc23858, nc23859, nc23860, 
        nc23861, nc23862, nc23863}), .DB_DETECT(\DB_DETECT[15][13] ), 
        .SB_CORRECT(\SB_CORRECT[15][13] ), .ACCESS_BUSY(
        \ACCESS_BUSY[15][13] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[27], W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C4 (.A_DOUT({nc23864, 
        nc23865, nc23866, nc23867, nc23868, nc23869, nc23870, nc23871, 
        nc23872, nc23873, nc23874, nc23875, nc23876, nc23877, nc23878, 
        nc23879, nc23880, nc23881, \R_DATA_TEMPR7[9] , 
        \R_DATA_TEMPR7[8] }), .B_DOUT({nc23882, nc23883, nc23884, 
        nc23885, nc23886, nc23887, nc23888, nc23889, nc23890, nc23891, 
        nc23892, nc23893, nc23894, nc23895, nc23896, nc23897, nc23898, 
        nc23899, nc23900, nc23901}), .DB_DETECT(\DB_DETECT[7][4] ), 
        .SB_CORRECT(\SB_CORRECT[7][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C7 (.A_DOUT({
        nc23902, nc23903, nc23904, nc23905, nc23906, nc23907, nc23908, 
        nc23909, nc23910, nc23911, nc23912, nc23913, nc23914, nc23915, 
        nc23916, nc23917, nc23918, nc23919, \R_DATA_TEMPR27[15] , 
        \R_DATA_TEMPR27[14] }), .B_DOUT({nc23920, nc23921, nc23922, 
        nc23923, nc23924, nc23925, nc23926, nc23927, nc23928, nc23929, 
        nc23930, nc23931, nc23932, nc23933, nc23934, nc23935, nc23936, 
        nc23937, nc23938, nc23939}), .DB_DETECT(\DB_DETECT[27][7] ), 
        .SB_CORRECT(\SB_CORRECT[27][7] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][7] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[15], W_DATA[14]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[7]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[28]  (.A(OR4_310_Y), .B(OR4_264_Y), .C(OR4_105_Y), 
        .D(OR4_143_Y), .Y(R_DATA[28]));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C12 (.A_DOUT({
        nc23940, nc23941, nc23942, nc23943, nc23944, nc23945, nc23946, 
        nc23947, nc23948, nc23949, nc23950, nc23951, nc23952, nc23953, 
        nc23954, nc23955, nc23956, nc23957, \R_DATA_TEMPR17[25] , 
        \R_DATA_TEMPR17[24] }), .B_DOUT({nc23958, nc23959, nc23960, 
        nc23961, nc23962, nc23963, nc23964, nc23965, nc23966, nc23967, 
        nc23968, nc23969, nc23970, nc23971, nc23972, nc23973, nc23974, 
        nc23975, nc23976, nc23977}), .DB_DETECT(\DB_DETECT[17][12] ), 
        .SB_CORRECT(\SB_CORRECT[17][12] ), .ACCESS_BUSY(
        \ACCESS_BUSY[17][12] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[25], W_DATA[24]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C11 (.A_DOUT({
        nc23978, nc23979, nc23980, nc23981, nc23982, nc23983, nc23984, 
        nc23985, nc23986, nc23987, nc23988, nc23989, nc23990, nc23991, 
        nc23992, nc23993, nc23994, nc23995, \R_DATA_TEMPR27[23] , 
        \R_DATA_TEMPR27[22] }), .B_DOUT({nc23996, nc23997, nc23998, 
        nc23999, nc24000, nc24001, nc24002, nc24003, nc24004, nc24005, 
        nc24006, nc24007, nc24008, nc24009, nc24010, nc24011, nc24012, 
        nc24013, nc24014, nc24015}), .DB_DETECT(\DB_DETECT[27][11] ), 
        .SB_CORRECT(\SB_CORRECT[27][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[27][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C17 (.A_DOUT({
        nc24016, nc24017, nc24018, nc24019, nc24020, nc24021, nc24022, 
        nc24023, nc24024, nc24025, nc24026, nc24027, nc24028, nc24029, 
        nc24030, nc24031, nc24032, nc24033, \R_DATA_TEMPR24[35] , 
        \R_DATA_TEMPR24[34] }), .B_DOUT({nc24034, nc24035, nc24036, 
        nc24037, nc24038, nc24039, nc24040, nc24041, nc24042, nc24043, 
        nc24044, nc24045, nc24046, nc24047, nc24048, nc24049, nc24050, 
        nc24051, nc24052, nc24053}), .DB_DETECT(\DB_DETECT[24][17] ), 
        .SB_CORRECT(\SB_CORRECT[24][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[24][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C3 (.A_DOUT({
        nc24054, nc24055, nc24056, nc24057, nc24058, nc24059, nc24060, 
        nc24061, nc24062, nc24063, nc24064, nc24065, nc24066, nc24067, 
        nc24068, nc24069, nc24070, nc24071, \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR21[6] }), .B_DOUT({nc24072, nc24073, nc24074, 
        nc24075, nc24076, nc24077, nc24078, nc24079, nc24080, nc24081, 
        nc24082, nc24083, nc24084, nc24085, nc24086, nc24087, nc24088, 
        nc24089, nc24090, nc24091}), .DB_DETECT(\DB_DETECT[21][3] ), 
        .SB_CORRECT(\SB_CORRECT[21][3] ), .ACCESS_BUSY(
        \ACCESS_BUSY[21][3] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[7], W_DATA[6]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C10 (.A_DOUT({
        nc24092, nc24093, nc24094, nc24095, nc24096, nc24097, nc24098, 
        nc24099, nc24100, nc24101, nc24102, nc24103, nc24104, nc24105, 
        nc24106, nc24107, nc24108, nc24109, \R_DATA_TEMPR4[21] , 
        \R_DATA_TEMPR4[20] }), .B_DOUT({nc24110, nc24111, nc24112, 
        nc24113, nc24114, nc24115, nc24116, nc24117, nc24118, nc24119, 
        nc24120, nc24121, nc24122, nc24123, nc24124, nc24125, nc24126, 
        nc24127, nc24128, nc24129}), .DB_DETECT(\DB_DETECT[4][10] ), 
        .SB_CORRECT(\SB_CORRECT[4][10] ), .ACCESS_BUSY(
        \ACCESS_BUSY[4][10] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[21], W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[10]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C11 (.A_DOUT({
        nc24130, nc24131, nc24132, nc24133, nc24134, nc24135, nc24136, 
        nc24137, nc24138, nc24139, nc24140, nc24141, nc24142, nc24143, 
        nc24144, nc24145, nc24146, nc24147, \R_DATA_TEMPR0[23] , 
        \R_DATA_TEMPR0[22] }), .B_DOUT({nc24148, nc24149, nc24150, 
        nc24151, nc24152, nc24153, nc24154, nc24155, nc24156, nc24157, 
        nc24158, nc24159, nc24160, nc24161, nc24162, nc24163, nc24164, 
        nc24165, nc24166, nc24167}), .DB_DETECT(\DB_DETECT[0][11] ), 
        .SB_CORRECT(\SB_CORRECT[0][11] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][11] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[0] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[23], W_DATA[22]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C8 (.A_DOUT({nc24168, 
        nc24169, nc24170, nc24171, nc24172, nc24173, nc24174, nc24175, 
        nc24176, nc24177, nc24178, nc24179, nc24180, nc24181, nc24182, 
        nc24183, nc24184, nc24185, \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR7[16] }), .B_DOUT({nc24186, nc24187, nc24188, 
        nc24189, nc24190, nc24191, nc24192, nc24193, nc24194, nc24195, 
        nc24196, nc24197, nc24198, nc24199, nc24200, nc24201, nc24202, 
        nc24203, nc24204, nc24205}), .DB_DETECT(\DB_DETECT[7][8] ), 
        .SB_CORRECT(\SB_CORRECT[7][8] ), .ACCESS_BUSY(
        \ACCESS_BUSY[7][8] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[1] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[17], W_DATA[16]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[8]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C17 (.A_DOUT({
        nc24206, nc24207, nc24208, nc24209, nc24210, nc24211, nc24212, 
        nc24213, nc24214, nc24215, nc24216, nc24217, nc24218, nc24219, 
        nc24220, nc24221, nc24222, nc24223, \R_DATA_TEMPR25[35] , 
        \R_DATA_TEMPR25[34] }), .B_DOUT({nc24224, nc24225, nc24226, 
        nc24227, nc24228, nc24229, nc24230, nc24231, nc24232, nc24233, 
        nc24234, nc24235, nc24236, nc24237, nc24238, nc24239, nc24240, 
        nc24241, nc24242, nc24243}), .DB_DETECT(\DB_DETECT[25][17] ), 
        .SB_CORRECT(\SB_CORRECT[25][17] ), .ACCESS_BUSY(
        \ACCESS_BUSY[25][17] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[35], W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_98 (.A(OR4_21_Y), .B(OR2_10_Y), .C(\R_DATA_TEMPR22[23] ), 
        .D(\R_DATA_TEMPR23[23] ), .Y(OR4_98_Y));
    OR4 OR4_321 (.A(\R_DATA_TEMPR28[31] ), .B(\R_DATA_TEMPR29[31] ), 
        .C(\R_DATA_TEMPR30[31] ), .D(\R_DATA_TEMPR31[31] ), .Y(
        OR4_321_Y));
    OR4 OR4_337 (.A(OR4_46_Y), .B(OR2_35_Y), .C(\R_DATA_TEMPR22[0] ), 
        .D(\R_DATA_TEMPR23[0] ), .Y(OR4_337_Y));
    OR4 OR4_130 (.A(OR4_53_Y), .B(OR2_38_Y), .C(\R_DATA_TEMPR22[13] ), 
        .D(\R_DATA_TEMPR23[13] ), .Y(OR4_130_Y));
    OR2 OR2_25 (.A(\R_DATA_TEMPR20[7] ), .B(\R_DATA_TEMPR21[7] ), .Y(
        OR2_25_Y));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C9 (.A_DOUT({
        nc24244, nc24245, nc24246, nc24247, nc24248, nc24249, nc24250, 
        nc24251, nc24252, nc24253, nc24254, nc24255, nc24256, nc24257, 
        nc24258, nc24259, nc24260, nc24261, \R_DATA_TEMPR14[19] , 
        \R_DATA_TEMPR14[18] }), .B_DOUT({nc24262, nc24263, nc24264, 
        nc24265, nc24266, nc24267, nc24268, nc24269, nc24270, nc24271, 
        nc24272, nc24273, nc24274, nc24275, nc24276, nc24277, nc24278, 
        nc24279, nc24280, nc24281}), .DB_DETECT(\DB_DETECT[14][9] ), 
        .SB_CORRECT(\SB_CORRECT[14][9] ), .ACCESS_BUSY(
        \ACCESS_BUSY[14][9] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[14], 
        \BLKY0[0] }), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[3] , 
        W_ADDR[14], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[19], W_DATA[18]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[9]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 lsram_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C4 (.A_DOUT({
        nc24282, nc24283, nc24284, nc24285, nc24286, nc24287, nc24288, 
        nc24289, nc24290, nc24291, nc24292, nc24293, nc24294, nc24295, 
        nc24296, nc24297, nc24298, nc24299, \R_DATA_TEMPR31[9] , 
        \R_DATA_TEMPR31[8] }), .B_DOUT({nc24300, nc24301, nc24302, 
        nc24303, nc24304, nc24305, nc24306, nc24307, nc24308, nc24309, 
        nc24310, nc24311, nc24312, nc24313, nc24314, nc24315, nc24316, 
        nc24317, nc24318, nc24319}), .DB_DETECT(\DB_DETECT[31][4] ), 
        .SB_CORRECT(\SB_CORRECT[31][4] ), .ACCESS_BUSY(
        \ACCESS_BUSY[31][4] ), .A_ADDR({R_ADDR[12], R_ADDR[11], 
        R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[14], 
        R_ADDR[13]}), .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .A_REN(VCC), .A_WEN({GND, GND}), .A_DOUT_EN(
        VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND}), .B_BLK_EN({\BLKX2[7] , 
        W_ADDR[14], W_ADDR[13]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, W_DATA[9], W_DATA[8]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[4]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_303 (.A(\R_DATA_TEMPR4[17] ), .B(\R_DATA_TEMPR5[17] ), .C(
        \R_DATA_TEMPR6[17] ), .D(\R_DATA_TEMPR7[17] ), .Y(OR4_303_Y));
    OR4 OR4_169 (.A(\R_DATA_TEMPR4[12] ), .B(\R_DATA_TEMPR5[12] ), .C(
        \R_DATA_TEMPR6[12] ), .D(\R_DATA_TEMPR7[12] ), .Y(OR4_169_Y));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
