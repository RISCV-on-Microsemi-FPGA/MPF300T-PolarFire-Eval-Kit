`timescale 1 ns/100 ps
// Version: PolarFire EAP4-SPA 12.100.8.13


module LSRAM_0_PF_URAM_0_PF_URAM(
       R_DATA,
       W_DATA,
       R_ADDR,
       W_ADDR,
       BLK_EN,
       CLK,
       W_EN
    );
output [39:0] R_DATA;
input  [39:0] W_DATA;
input  [10:0] R_ADDR;
input  [10:0] W_ADDR;
input  BLK_EN;
input  CLK;
input  W_EN;

    wire \R_DATA_TEMPR0[0] , \R_DATA_TEMPR1[0] , \R_DATA_TEMPR2[0] , 
        \R_DATA_TEMPR3[0] , \R_DATA_TEMPR4[0] , \R_DATA_TEMPR5[0] , 
        \R_DATA_TEMPR6[0] , \R_DATA_TEMPR7[0] , \R_DATA_TEMPR8[0] , 
        \R_DATA_TEMPR9[0] , \R_DATA_TEMPR10[0] , \R_DATA_TEMPR11[0] , 
        \R_DATA_TEMPR12[0] , \R_DATA_TEMPR13[0] , \R_DATA_TEMPR14[0] , 
        \R_DATA_TEMPR15[0] , \R_DATA_TEMPR16[0] , \R_DATA_TEMPR17[0] , 
        \R_DATA_TEMPR18[0] , \R_DATA_TEMPR19[0] , \R_DATA_TEMPR20[0] , 
        \R_DATA_TEMPR21[0] , \R_DATA_TEMPR22[0] , \R_DATA_TEMPR23[0] , 
        \R_DATA_TEMPR24[0] , \R_DATA_TEMPR25[0] , \R_DATA_TEMPR26[0] , 
        \R_DATA_TEMPR27[0] , \R_DATA_TEMPR28[0] , \R_DATA_TEMPR29[0] , 
        \R_DATA_TEMPR30[0] , \R_DATA_TEMPR31[0] , \R_DATA_TEMPR0[1] , 
        \R_DATA_TEMPR1[1] , \R_DATA_TEMPR2[1] , \R_DATA_TEMPR3[1] , 
        \R_DATA_TEMPR4[1] , \R_DATA_TEMPR5[1] , \R_DATA_TEMPR6[1] , 
        \R_DATA_TEMPR7[1] , \R_DATA_TEMPR8[1] , \R_DATA_TEMPR9[1] , 
        \R_DATA_TEMPR10[1] , \R_DATA_TEMPR11[1] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR13[1] , \R_DATA_TEMPR14[1] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR16[1] , \R_DATA_TEMPR17[1] , \R_DATA_TEMPR18[1] , 
        \R_DATA_TEMPR19[1] , \R_DATA_TEMPR20[1] , \R_DATA_TEMPR21[1] , 
        \R_DATA_TEMPR22[1] , \R_DATA_TEMPR23[1] , \R_DATA_TEMPR24[1] , 
        \R_DATA_TEMPR25[1] , \R_DATA_TEMPR26[1] , \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR28[1] , \R_DATA_TEMPR29[1] , \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR31[1] , \R_DATA_TEMPR0[2] , \R_DATA_TEMPR1[2] , 
        \R_DATA_TEMPR2[2] , \R_DATA_TEMPR3[2] , \R_DATA_TEMPR4[2] , 
        \R_DATA_TEMPR5[2] , \R_DATA_TEMPR6[2] , \R_DATA_TEMPR7[2] , 
        \R_DATA_TEMPR8[2] , \R_DATA_TEMPR9[2] , \R_DATA_TEMPR10[2] , 
        \R_DATA_TEMPR11[2] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR13[2] , 
        \R_DATA_TEMPR14[2] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR16[2] , 
        \R_DATA_TEMPR17[2] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR19[2] , 
        \R_DATA_TEMPR20[2] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR22[2] , 
        \R_DATA_TEMPR23[2] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR25[2] , 
        \R_DATA_TEMPR26[2] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR28[2] , 
        \R_DATA_TEMPR29[2] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR31[2] , 
        \R_DATA_TEMPR0[3] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR2[3] , 
        \R_DATA_TEMPR3[3] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR5[3] , 
        \R_DATA_TEMPR6[3] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR8[3] , 
        \R_DATA_TEMPR9[3] , \R_DATA_TEMPR10[3] , \R_DATA_TEMPR11[3] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR13[3] , \R_DATA_TEMPR14[3] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR16[3] , \R_DATA_TEMPR17[3] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR19[3] , \R_DATA_TEMPR20[3] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR22[3] , \R_DATA_TEMPR23[3] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR25[3] , \R_DATA_TEMPR26[3] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR28[3] , \R_DATA_TEMPR29[3] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR31[3] , \R_DATA_TEMPR0[4] , 
        \R_DATA_TEMPR1[4] , \R_DATA_TEMPR2[4] , \R_DATA_TEMPR3[4] , 
        \R_DATA_TEMPR4[4] , \R_DATA_TEMPR5[4] , \R_DATA_TEMPR6[4] , 
        \R_DATA_TEMPR7[4] , \R_DATA_TEMPR8[4] , \R_DATA_TEMPR9[4] , 
        \R_DATA_TEMPR10[4] , \R_DATA_TEMPR11[4] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR13[4] , \R_DATA_TEMPR14[4] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR16[4] , \R_DATA_TEMPR17[4] , \R_DATA_TEMPR18[4] , 
        \R_DATA_TEMPR19[4] , \R_DATA_TEMPR20[4] , \R_DATA_TEMPR21[4] , 
        \R_DATA_TEMPR22[4] , \R_DATA_TEMPR23[4] , \R_DATA_TEMPR24[4] , 
        \R_DATA_TEMPR25[4] , \R_DATA_TEMPR26[4] , \R_DATA_TEMPR27[4] , 
        \R_DATA_TEMPR28[4] , \R_DATA_TEMPR29[4] , \R_DATA_TEMPR30[4] , 
        \R_DATA_TEMPR31[4] , \R_DATA_TEMPR0[5] , \R_DATA_TEMPR1[5] , 
        \R_DATA_TEMPR2[5] , \R_DATA_TEMPR3[5] , \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR5[5] , \R_DATA_TEMPR6[5] , \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR8[5] , \R_DATA_TEMPR9[5] , \R_DATA_TEMPR10[5] , 
        \R_DATA_TEMPR11[5] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR13[5] , 
        \R_DATA_TEMPR14[5] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR16[5] , 
        \R_DATA_TEMPR17[5] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR19[5] , 
        \R_DATA_TEMPR20[5] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR22[5] , 
        \R_DATA_TEMPR23[5] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR25[5] , 
        \R_DATA_TEMPR26[5] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR28[5] , 
        \R_DATA_TEMPR29[5] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR31[5] , 
        \R_DATA_TEMPR0[6] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR2[6] , 
        \R_DATA_TEMPR3[6] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR5[6] , 
        \R_DATA_TEMPR6[6] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR8[6] , 
        \R_DATA_TEMPR9[6] , \R_DATA_TEMPR10[6] , \R_DATA_TEMPR11[6] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR13[6] , \R_DATA_TEMPR14[6] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR16[6] , \R_DATA_TEMPR17[6] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR19[6] , \R_DATA_TEMPR20[6] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR22[6] , \R_DATA_TEMPR23[6] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR25[6] , \R_DATA_TEMPR26[6] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR28[6] , \R_DATA_TEMPR29[6] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR31[6] , \R_DATA_TEMPR0[7] , 
        \R_DATA_TEMPR1[7] , \R_DATA_TEMPR2[7] , \R_DATA_TEMPR3[7] , 
        \R_DATA_TEMPR4[7] , \R_DATA_TEMPR5[7] , \R_DATA_TEMPR6[7] , 
        \R_DATA_TEMPR7[7] , \R_DATA_TEMPR8[7] , \R_DATA_TEMPR9[7] , 
        \R_DATA_TEMPR10[7] , \R_DATA_TEMPR11[7] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR13[7] , \R_DATA_TEMPR14[7] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR16[7] , \R_DATA_TEMPR17[7] , \R_DATA_TEMPR18[7] , 
        \R_DATA_TEMPR19[7] , \R_DATA_TEMPR20[7] , \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR22[7] , \R_DATA_TEMPR23[7] , \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR25[7] , \R_DATA_TEMPR26[7] , \R_DATA_TEMPR27[7] , 
        \R_DATA_TEMPR28[7] , \R_DATA_TEMPR29[7] , \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR31[7] , \R_DATA_TEMPR0[8] , \R_DATA_TEMPR1[8] , 
        \R_DATA_TEMPR2[8] , \R_DATA_TEMPR3[8] , \R_DATA_TEMPR4[8] , 
        \R_DATA_TEMPR5[8] , \R_DATA_TEMPR6[8] , \R_DATA_TEMPR7[8] , 
        \R_DATA_TEMPR8[8] , \R_DATA_TEMPR9[8] , \R_DATA_TEMPR10[8] , 
        \R_DATA_TEMPR11[8] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR13[8] , 
        \R_DATA_TEMPR14[8] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR16[8] , 
        \R_DATA_TEMPR17[8] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR19[8] , 
        \R_DATA_TEMPR20[8] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR22[8] , 
        \R_DATA_TEMPR23[8] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR25[8] , 
        \R_DATA_TEMPR26[8] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR28[8] , 
        \R_DATA_TEMPR29[8] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR31[8] , 
        \R_DATA_TEMPR0[9] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR2[9] , 
        \R_DATA_TEMPR3[9] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR5[9] , 
        \R_DATA_TEMPR6[9] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR8[9] , 
        \R_DATA_TEMPR9[9] , \R_DATA_TEMPR10[9] , \R_DATA_TEMPR11[9] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR13[9] , \R_DATA_TEMPR14[9] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR16[9] , \R_DATA_TEMPR17[9] , 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR19[9] , \R_DATA_TEMPR20[9] , 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR22[9] , \R_DATA_TEMPR23[9] , 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR25[9] , \R_DATA_TEMPR26[9] , 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR28[9] , \R_DATA_TEMPR29[9] , 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR31[9] , \R_DATA_TEMPR0[10] , 
        \R_DATA_TEMPR1[10] , \R_DATA_TEMPR2[10] , \R_DATA_TEMPR3[10] , 
        \R_DATA_TEMPR4[10] , \R_DATA_TEMPR5[10] , \R_DATA_TEMPR6[10] , 
        \R_DATA_TEMPR7[10] , \R_DATA_TEMPR8[10] , \R_DATA_TEMPR9[10] , 
        \R_DATA_TEMPR10[10] , \R_DATA_TEMPR11[10] , 
        \R_DATA_TEMPR12[10] , \R_DATA_TEMPR13[10] , 
        \R_DATA_TEMPR14[10] , \R_DATA_TEMPR15[10] , 
        \R_DATA_TEMPR16[10] , \R_DATA_TEMPR17[10] , 
        \R_DATA_TEMPR18[10] , \R_DATA_TEMPR19[10] , 
        \R_DATA_TEMPR20[10] , \R_DATA_TEMPR21[10] , 
        \R_DATA_TEMPR22[10] , \R_DATA_TEMPR23[10] , 
        \R_DATA_TEMPR24[10] , \R_DATA_TEMPR25[10] , 
        \R_DATA_TEMPR26[10] , \R_DATA_TEMPR27[10] , 
        \R_DATA_TEMPR28[10] , \R_DATA_TEMPR29[10] , 
        \R_DATA_TEMPR30[10] , \R_DATA_TEMPR31[10] , 
        \R_DATA_TEMPR0[11] , \R_DATA_TEMPR1[11] , \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR3[11] , \R_DATA_TEMPR4[11] , \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR6[11] , \R_DATA_TEMPR7[11] , \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR9[11] , \R_DATA_TEMPR10[11] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR12[11] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR14[11] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR16[11] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR18[11] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR20[11] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR22[11] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR24[11] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR26[11] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR28[11] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR30[11] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR1[12] , 
        \R_DATA_TEMPR2[12] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR4[12] , 
        \R_DATA_TEMPR5[12] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR7[12] , 
        \R_DATA_TEMPR8[12] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR11[12] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR13[12] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR15[12] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR17[12] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR19[12] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR21[12] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR23[12] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR25[12] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR27[12] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR29[12] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR31[12] , \R_DATA_TEMPR0[13] , \R_DATA_TEMPR1[13] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR3[13] , \R_DATA_TEMPR4[13] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR6[13] , \R_DATA_TEMPR7[13] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR9[13] , \R_DATA_TEMPR10[13] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR12[13] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR14[13] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR16[13] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR18[13] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR20[13] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR22[13] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR24[13] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR26[13] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR28[13] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR30[13] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR0[14] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR2[14] , \R_DATA_TEMPR3[14] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR5[14] , \R_DATA_TEMPR6[14] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR8[14] , \R_DATA_TEMPR9[14] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR11[14] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR13[14] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR15[14] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR17[14] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR19[14] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR21[14] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR23[14] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR25[14] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR27[14] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR29[14] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR31[14] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR1[15] , 
        \R_DATA_TEMPR2[15] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR4[15] , 
        \R_DATA_TEMPR5[15] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR7[15] , 
        \R_DATA_TEMPR8[15] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR10[15] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR12[15] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR14[15] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR16[15] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR18[15] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR20[15] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR22[15] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR24[15] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR26[15] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR28[15] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR30[15] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR0[16] , \R_DATA_TEMPR1[16] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR3[16] , \R_DATA_TEMPR4[16] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR6[16] , \R_DATA_TEMPR7[16] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR9[16] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR11[16] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR13[16] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR15[16] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR17[16] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR19[16] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR21[16] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR23[16] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR25[16] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR27[16] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR29[16] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR31[16] , \R_DATA_TEMPR0[17] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR2[17] , \R_DATA_TEMPR3[17] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR5[17] , \R_DATA_TEMPR6[17] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR8[17] , \R_DATA_TEMPR9[17] , \R_DATA_TEMPR10[17] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR12[17] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR14[17] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR16[17] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR18[17] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR20[17] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR22[17] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR24[17] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR26[17] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR28[17] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR30[17] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR1[18] , 
        \R_DATA_TEMPR2[18] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR4[18] , 
        \R_DATA_TEMPR5[18] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR7[18] , 
        \R_DATA_TEMPR8[18] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR11[18] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR13[18] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR15[18] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR17[18] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR19[18] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR21[18] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR23[18] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR25[18] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR27[18] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR29[18] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR31[18] , \R_DATA_TEMPR0[19] , \R_DATA_TEMPR1[19] , 
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR3[19] , \R_DATA_TEMPR4[19] , 
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR6[19] , \R_DATA_TEMPR7[19] , 
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR9[19] , \R_DATA_TEMPR10[19] , 
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR12[19] , 
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR14[19] , 
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR16[19] , 
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR18[19] , 
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR20[19] , 
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR22[19] , 
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR24[19] , 
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR26[19] , 
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR28[19] , 
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR30[19] , 
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR0[20] , \R_DATA_TEMPR1[20] , 
        \R_DATA_TEMPR2[20] , \R_DATA_TEMPR3[20] , \R_DATA_TEMPR4[20] , 
        \R_DATA_TEMPR5[20] , \R_DATA_TEMPR6[20] , \R_DATA_TEMPR7[20] , 
        \R_DATA_TEMPR8[20] , \R_DATA_TEMPR9[20] , \R_DATA_TEMPR10[20] , 
        \R_DATA_TEMPR11[20] , \R_DATA_TEMPR12[20] , 
        \R_DATA_TEMPR13[20] , \R_DATA_TEMPR14[20] , 
        \R_DATA_TEMPR15[20] , \R_DATA_TEMPR16[20] , 
        \R_DATA_TEMPR17[20] , \R_DATA_TEMPR18[20] , 
        \R_DATA_TEMPR19[20] , \R_DATA_TEMPR20[20] , 
        \R_DATA_TEMPR21[20] , \R_DATA_TEMPR22[20] , 
        \R_DATA_TEMPR23[20] , \R_DATA_TEMPR24[20] , 
        \R_DATA_TEMPR25[20] , \R_DATA_TEMPR26[20] , 
        \R_DATA_TEMPR27[20] , \R_DATA_TEMPR28[20] , 
        \R_DATA_TEMPR29[20] , \R_DATA_TEMPR30[20] , 
        \R_DATA_TEMPR31[20] , \R_DATA_TEMPR0[21] , \R_DATA_TEMPR1[21] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR3[21] , \R_DATA_TEMPR4[21] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR6[21] , \R_DATA_TEMPR7[21] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR9[21] , \R_DATA_TEMPR10[21] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR12[21] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR14[21] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR16[21] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR18[21] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR20[21] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR22[21] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR24[21] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR26[21] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR28[21] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR30[21] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR0[22] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR2[22] , \R_DATA_TEMPR3[22] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR5[22] , \R_DATA_TEMPR6[22] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR8[22] , \R_DATA_TEMPR9[22] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR11[22] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR13[22] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR15[22] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR17[22] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR19[22] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR21[22] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR23[22] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR25[22] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR27[22] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR29[22] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR31[22] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR1[23] , 
        \R_DATA_TEMPR2[23] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR4[23] , 
        \R_DATA_TEMPR5[23] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR7[23] , 
        \R_DATA_TEMPR8[23] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR10[23] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR12[23] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR14[23] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR16[23] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR18[23] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR20[23] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR22[23] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR24[23] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR26[23] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR28[23] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR30[23] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR0[24] , \R_DATA_TEMPR1[24] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR3[24] , \R_DATA_TEMPR4[24] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR6[24] , \R_DATA_TEMPR7[24] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR9[24] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR11[24] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR13[24] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR15[24] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR17[24] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR19[24] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR21[24] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR23[24] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR25[24] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR27[24] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR29[24] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR31[24] , \R_DATA_TEMPR0[25] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR2[25] , \R_DATA_TEMPR3[25] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR5[25] , \R_DATA_TEMPR6[25] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR8[25] , \R_DATA_TEMPR9[25] , \R_DATA_TEMPR10[25] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR12[25] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR14[25] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR16[25] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR18[25] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR20[25] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR22[25] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR24[25] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR26[25] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR28[25] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR30[25] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR1[26] , 
        \R_DATA_TEMPR2[26] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR4[26] , 
        \R_DATA_TEMPR5[26] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR7[26] , 
        \R_DATA_TEMPR8[26] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR11[26] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR13[26] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR15[26] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR17[26] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR19[26] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR21[26] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR23[26] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR25[26] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR27[26] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR29[26] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR31[26] , \R_DATA_TEMPR0[27] , \R_DATA_TEMPR1[27] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR3[27] , \R_DATA_TEMPR4[27] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR6[27] , \R_DATA_TEMPR7[27] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR9[27] , \R_DATA_TEMPR10[27] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR12[27] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR14[27] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR16[27] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR18[27] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR20[27] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR22[27] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR24[27] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR26[27] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR28[27] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR30[27] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR0[28] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR2[28] , \R_DATA_TEMPR3[28] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR5[28] , \R_DATA_TEMPR6[28] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR8[28] , \R_DATA_TEMPR9[28] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR11[28] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR13[28] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR15[28] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR17[28] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR19[28] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR21[28] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR23[28] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR25[28] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR27[28] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR29[28] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR31[28] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR1[29] , 
        \R_DATA_TEMPR2[29] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR4[29] , 
        \R_DATA_TEMPR5[29] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR7[29] , 
        \R_DATA_TEMPR8[29] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR10[29] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR12[29] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR14[29] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR16[29] , 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR18[29] , 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR20[29] , 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR22[29] , 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR24[29] , 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR26[29] , 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR28[29] , 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR30[29] , 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR0[30] , \R_DATA_TEMPR1[30] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR3[30] , \R_DATA_TEMPR4[30] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR6[30] , \R_DATA_TEMPR7[30] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR9[30] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR11[30] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR13[30] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR15[30] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR17[30] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR19[30] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR21[30] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR23[30] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR25[30] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR27[30] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR29[30] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR31[30] , \R_DATA_TEMPR0[31] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR2[31] , \R_DATA_TEMPR3[31] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR5[31] , \R_DATA_TEMPR6[31] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR8[31] , \R_DATA_TEMPR9[31] , \R_DATA_TEMPR10[31] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR12[31] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR14[31] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR16[31] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR18[31] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR20[31] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR22[31] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR24[31] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR26[31] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR28[31] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR30[31] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR1[32] , 
        \R_DATA_TEMPR2[32] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR4[32] , 
        \R_DATA_TEMPR5[32] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR7[32] , 
        \R_DATA_TEMPR8[32] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR11[32] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR13[32] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR15[32] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR17[32] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR19[32] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR21[32] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR23[32] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR25[32] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR27[32] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR29[32] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR31[32] , \R_DATA_TEMPR0[33] , \R_DATA_TEMPR1[33] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR3[33] , \R_DATA_TEMPR4[33] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR6[33] , \R_DATA_TEMPR7[33] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR9[33] , \R_DATA_TEMPR10[33] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR12[33] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR14[33] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR16[33] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR18[33] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR20[33] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR22[33] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR24[33] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR26[33] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR28[33] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR30[33] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR0[34] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR2[34] , \R_DATA_TEMPR3[34] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR5[34] , \R_DATA_TEMPR6[34] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR8[34] , \R_DATA_TEMPR9[34] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR11[34] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR13[34] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR15[34] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR17[34] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR19[34] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR21[34] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR23[34] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR25[34] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR27[34] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR29[34] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR31[34] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR1[35] , 
        \R_DATA_TEMPR2[35] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR4[35] , 
        \R_DATA_TEMPR5[35] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR7[35] , 
        \R_DATA_TEMPR8[35] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR10[35] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR12[35] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR14[35] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR16[35] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR18[35] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR20[35] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR22[35] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR24[35] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR26[35] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR28[35] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR30[35] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR0[36] , \R_DATA_TEMPR1[36] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR3[36] , \R_DATA_TEMPR4[36] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR6[36] , \R_DATA_TEMPR7[36] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR9[36] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR11[36] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR13[36] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR15[36] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR17[36] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR19[36] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR21[36] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR23[36] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR25[36] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR27[36] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR29[36] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR31[36] , \R_DATA_TEMPR0[37] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR2[37] , \R_DATA_TEMPR3[37] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR5[37] , \R_DATA_TEMPR6[37] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR8[37] , \R_DATA_TEMPR9[37] , \R_DATA_TEMPR10[37] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR12[37] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR14[37] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR16[37] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR18[37] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR20[37] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR22[37] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR24[37] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR26[37] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR28[37] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR30[37] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR1[38] , 
        \R_DATA_TEMPR2[38] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR4[38] , 
        \R_DATA_TEMPR5[38] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR7[38] , 
        \R_DATA_TEMPR8[38] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR11[38] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR13[38] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR15[38] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR17[38] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR19[38] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR21[38] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR23[38] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR25[38] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR27[38] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR29[38] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR31[38] , \R_DATA_TEMPR0[39] , \R_DATA_TEMPR1[39] , 
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR3[39] , \R_DATA_TEMPR4[39] , 
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR6[39] , \R_DATA_TEMPR7[39] , 
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR9[39] , \R_DATA_TEMPR10[39] , 
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR12[39] , 
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR14[39] , 
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR16[39] , 
        \R_DATA_TEMPR17[39] , \R_DATA_TEMPR18[39] , 
        \R_DATA_TEMPR19[39] , \R_DATA_TEMPR20[39] , 
        \R_DATA_TEMPR21[39] , \R_DATA_TEMPR22[39] , 
        \R_DATA_TEMPR23[39] , \R_DATA_TEMPR24[39] , 
        \R_DATA_TEMPR25[39] , \R_DATA_TEMPR26[39] , 
        \R_DATA_TEMPR27[39] , \R_DATA_TEMPR28[39] , 
        \R_DATA_TEMPR29[39] , \R_DATA_TEMPR30[39] , 
        \R_DATA_TEMPR31[39] , \BLKX0[0] , \BLKX0[1] , \BLKX0[2] , 
        \BLKX0[3] , \BLKX0[4] , \BLKX0[5] , \BLKX0[6] , \BLKX0[7] , 
        \BLKX0[8] , \BLKX0[9] , \BLKX0[10] , \BLKX0[11] , \BLKX0[12] , 
        \BLKX0[13] , \BLKX0[14] , \BLKX0[15] , \BLKX0[16] , 
        \BLKX0[17] , \BLKX0[18] , \BLKX0[19] , \BLKX0[20] , 
        \BLKX0[21] , \BLKX0[22] , \BLKX0[23] , \BLKX0[24] , 
        \BLKX0[25] , \BLKX0[26] , \BLKX0[27] , \BLKX0[28] , 
        \BLKX0[29] , \BLKX0[30] , \BLKX0[31] , \BLKZ0[0] , \BLKZ0[1] , 
        \BLKZ0[2] , \BLKZ0[3] , \BLKZ0[4] , \BLKZ0[5] , \BLKZ0[6] , 
        \BLKZ0[7] , \BLKZ0[8] , \BLKZ0[9] , \BLKZ0[10] , \BLKZ0[11] , 
        \BLKZ0[12] , \BLKZ0[13] , \BLKZ0[14] , \BLKZ0[15] , 
        \BLKZ0[16] , \BLKZ0[17] , \BLKZ0[18] , \BLKZ0[19] , 
        \BLKZ0[20] , \BLKZ0[21] , \BLKZ0[22] , \BLKZ0[23] , 
        \BLKZ0[24] , \BLKZ0[25] , \BLKZ0[26] , \BLKZ0[27] , 
        \BLKZ0[28] , \BLKZ0[29] , \BLKZ0[30] , \BLKZ0[31] , 
        \ACCESS_BUSY[0][0] , \ACCESS_BUSY[0][1] , \ACCESS_BUSY[0][2] , 
        \ACCESS_BUSY[0][3] , \ACCESS_BUSY[1][0] , \ACCESS_BUSY[1][1] , 
        \ACCESS_BUSY[1][2] , \ACCESS_BUSY[1][3] , \ACCESS_BUSY[2][0] , 
        \ACCESS_BUSY[2][1] , \ACCESS_BUSY[2][2] , \ACCESS_BUSY[2][3] , 
        \ACCESS_BUSY[3][0] , \ACCESS_BUSY[3][1] , \ACCESS_BUSY[3][2] , 
        \ACCESS_BUSY[3][3] , \ACCESS_BUSY[4][0] , \ACCESS_BUSY[4][1] , 
        \ACCESS_BUSY[4][2] , \ACCESS_BUSY[4][3] , \ACCESS_BUSY[5][0] , 
        \ACCESS_BUSY[5][1] , \ACCESS_BUSY[5][2] , \ACCESS_BUSY[5][3] , 
        \ACCESS_BUSY[6][0] , \ACCESS_BUSY[6][1] , \ACCESS_BUSY[6][2] , 
        \ACCESS_BUSY[6][3] , \ACCESS_BUSY[7][0] , \ACCESS_BUSY[7][1] , 
        \ACCESS_BUSY[7][2] , \ACCESS_BUSY[7][3] , \ACCESS_BUSY[8][0] , 
        \ACCESS_BUSY[8][1] , \ACCESS_BUSY[8][2] , \ACCESS_BUSY[8][3] , 
        \ACCESS_BUSY[9][0] , \ACCESS_BUSY[9][1] , \ACCESS_BUSY[9][2] , 
        \ACCESS_BUSY[9][3] , \ACCESS_BUSY[10][0] , 
        \ACCESS_BUSY[10][1] , \ACCESS_BUSY[10][2] , 
        \ACCESS_BUSY[10][3] , \ACCESS_BUSY[11][0] , 
        \ACCESS_BUSY[11][1] , \ACCESS_BUSY[11][2] , 
        \ACCESS_BUSY[11][3] , \ACCESS_BUSY[12][0] , 
        \ACCESS_BUSY[12][1] , \ACCESS_BUSY[12][2] , 
        \ACCESS_BUSY[12][3] , \ACCESS_BUSY[13][0] , 
        \ACCESS_BUSY[13][1] , \ACCESS_BUSY[13][2] , 
        \ACCESS_BUSY[13][3] , \ACCESS_BUSY[14][0] , 
        \ACCESS_BUSY[14][1] , \ACCESS_BUSY[14][2] , 
        \ACCESS_BUSY[14][3] , \ACCESS_BUSY[15][0] , 
        \ACCESS_BUSY[15][1] , \ACCESS_BUSY[15][2] , 
        \ACCESS_BUSY[15][3] , \ACCESS_BUSY[16][0] , 
        \ACCESS_BUSY[16][1] , \ACCESS_BUSY[16][2] , 
        \ACCESS_BUSY[16][3] , \ACCESS_BUSY[17][0] , 
        \ACCESS_BUSY[17][1] , \ACCESS_BUSY[17][2] , 
        \ACCESS_BUSY[17][3] , \ACCESS_BUSY[18][0] , 
        \ACCESS_BUSY[18][1] , \ACCESS_BUSY[18][2] , 
        \ACCESS_BUSY[18][3] , \ACCESS_BUSY[19][0] , 
        \ACCESS_BUSY[19][1] , \ACCESS_BUSY[19][2] , 
        \ACCESS_BUSY[19][3] , \ACCESS_BUSY[20][0] , 
        \ACCESS_BUSY[20][1] , \ACCESS_BUSY[20][2] , 
        \ACCESS_BUSY[20][3] , \ACCESS_BUSY[21][0] , 
        \ACCESS_BUSY[21][1] , \ACCESS_BUSY[21][2] , 
        \ACCESS_BUSY[21][3] , \ACCESS_BUSY[22][0] , 
        \ACCESS_BUSY[22][1] , \ACCESS_BUSY[22][2] , 
        \ACCESS_BUSY[22][3] , \ACCESS_BUSY[23][0] , 
        \ACCESS_BUSY[23][1] , \ACCESS_BUSY[23][2] , 
        \ACCESS_BUSY[23][3] , \ACCESS_BUSY[24][0] , 
        \ACCESS_BUSY[24][1] , \ACCESS_BUSY[24][2] , 
        \ACCESS_BUSY[24][3] , \ACCESS_BUSY[25][0] , 
        \ACCESS_BUSY[25][1] , \ACCESS_BUSY[25][2] , 
        \ACCESS_BUSY[25][3] , \ACCESS_BUSY[26][0] , 
        \ACCESS_BUSY[26][1] , \ACCESS_BUSY[26][2] , 
        \ACCESS_BUSY[26][3] , \ACCESS_BUSY[27][0] , 
        \ACCESS_BUSY[27][1] , \ACCESS_BUSY[27][2] , 
        \ACCESS_BUSY[27][3] , \ACCESS_BUSY[28][0] , 
        \ACCESS_BUSY[28][1] , \ACCESS_BUSY[28][2] , 
        \ACCESS_BUSY[28][3] , \ACCESS_BUSY[29][0] , 
        \ACCESS_BUSY[29][1] , \ACCESS_BUSY[29][2] , 
        \ACCESS_BUSY[29][3] , \ACCESS_BUSY[30][0] , 
        \ACCESS_BUSY[30][1] , \ACCESS_BUSY[30][2] , 
        \ACCESS_BUSY[30][3] , \ACCESS_BUSY[31][0] , 
        \ACCESS_BUSY[31][1] , \ACCESS_BUSY[31][2] , 
        \ACCESS_BUSY[31][3] , OR4_192_Y, OR4_170_Y, OR4_243_Y, 
        OR4_274_Y, OR4_231_Y, OR4_113_Y, OR4_234_Y, OR4_104_Y, 
        OR4_240_Y, OR2_23_Y, OR4_40_Y, OR4_211_Y, OR4_306_Y, OR4_347_Y, 
        OR4_76_Y, OR4_276_Y, OR4_45_Y, OR4_219_Y, OR4_161_Y, OR2_36_Y, 
        OR4_14_Y, OR4_103_Y, OR4_259_Y, OR4_128_Y, OR4_354_Y, 
        OR4_272_Y, OR4_358_Y, OR4_148_Y, OR4_144_Y, OR2_11_Y, 
        OR4_301_Y, OR4_205_Y, OR4_191_Y, OR4_176_Y, OR4_54_Y, 
        OR4_357_Y, OR4_348_Y, OR4_200_Y, OR4_137_Y, OR2_1_Y, OR4_89_Y, 
        OR4_180_Y, OR4_151_Y, OR4_179_Y, OR4_110_Y, OR4_221_Y, 
        OR4_316_Y, OR4_123_Y, OR4_139_Y, OR2_9_Y, OR4_60_Y, OR4_15_Y, 
        OR4_208_Y, OR4_260_Y, OR4_314_Y, OR4_239_Y, OR4_175_Y, 
        OR4_194_Y, OR4_183_Y, OR2_18_Y, OR4_174_Y, OR4_214_Y, 
        OR4_134_Y, OR4_269_Y, OR4_47_Y, OR4_75_Y, OR4_190_Y, OR4_71_Y, 
        OR4_235_Y, OR2_21_Y, OR4_135_Y, OR4_331_Y, OR4_28_Y, OR4_48_Y, 
        OR4_307_Y, OR4_199_Y, OR4_217_Y, OR4_289_Y, OR4_49_Y, OR2_2_Y, 
        OR4_84_Y, OR4_3_Y, OR4_338_Y, OR4_280_Y, OR4_223_Y, OR4_355_Y, 
        OR4_138_Y, OR4_291_Y, OR4_155_Y, OR2_39_Y, OR4_51_Y, OR4_343_Y, 
        OR4_222_Y, OR4_298_Y, OR4_157_Y, OR4_288_Y, OR4_252_Y, 
        OR4_112_Y, OR4_50_Y, OR2_5_Y, OR4_83_Y, OR4_61_Y, OR4_70_Y, 
        OR4_321_Y, OR4_201_Y, OR4_267_Y, OR4_265_Y, OR4_323_Y, 
        OR4_165_Y, OR2_19_Y, OR4_225_Y, OR4_213_Y, OR4_163_Y, OR4_7_Y, 
        OR4_296_Y, OR4_140_Y, OR4_216_Y, OR4_36_Y, OR4_62_Y, OR2_16_Y, 
        OR4_77_Y, OR4_244_Y, OR4_339_Y, OR4_12_Y, OR4_109_Y, OR4_303_Y, 
        OR4_81_Y, OR4_250_Y, OR4_195_Y, OR2_24_Y, OR4_285_Y, OR4_97_Y, 
        OR4_230_Y, OR4_133_Y, OR4_59_Y, OR4_275_Y, OR4_290_Y, 
        OR4_115_Y, OR4_313_Y, OR2_22_Y, OR4_206_Y, OR4_325_Y, 
        OR4_224_Y, OR4_167_Y, OR4_350_Y, OR4_44_Y, OR4_261_Y, 
        OR4_215_Y, OR4_101_Y, OR2_25_Y, OR4_160_Y, OR4_2_Y, OR4_63_Y, 
        OR4_86_Y, OR4_340_Y, OR4_229_Y, OR4_248_Y, OR4_318_Y, OR4_91_Y, 
        OR2_33_Y, OR4_117_Y, OR4_26_Y, OR4_9_Y, OR4_304_Y, OR4_254_Y, 
        OR4_16_Y, OR4_166_Y, OR4_322_Y, OR4_189_Y, OR2_28_Y, OR4_292_Y, 
        OR4_334_Y, OR4_236_Y, OR4_188_Y, OR4_326_Y, OR4_4_Y, OR4_24_Y, 
        OR4_6_Y, OR4_209_Y, OR2_34_Y, OR4_256_Y, OR4_245_Y, OR4_196_Y, 
        OR4_29_Y, OR4_324_Y, OR4_169_Y, OR4_247_Y, OR4_72_Y, OR4_100_Y, 
        OR2_0_Y, OR4_312_Y, OR4_129_Y, OR4_263_Y, OR4_156_Y, OR4_96_Y, 
        OR4_302_Y, OR4_319_Y, OR4_136_Y, OR4_349_Y, OR2_7_Y, OR4_308_Y, 
        OR4_181_Y, OR4_1_Y, OR4_152_Y, OR4_249_Y, OR4_327_Y, OR4_8_Y, 
        OR4_273_Y, OR4_284_Y, OR2_26_Y, OR4_41_Y, OR4_118_Y, OR4_203_Y, 
        OR4_279_Y, OR4_116_Y, OR4_315_Y, OR4_197_Y, OR4_78_Y, 
        OR4_182_Y, OR2_3_Y, OR4_153_Y, OR4_329_Y, OR4_56_Y, OR4_99_Y, 
        OR4_184_Y, OR4_19_Y, OR4_159_Y, OR4_335_Y, OR4_281_Y, OR2_30_Y, 
        OR4_297_Y, OR4_337_Y, OR4_220_Y, OR4_293_Y, OR4_287_Y, 
        OR4_283_Y, OR4_255_Y, OR4_353_Y, OR4_46_Y, OR2_35_Y, OR4_262_Y, 
        OR4_351_Y, OR4_141_Y, OR4_10_Y, OR4_232_Y, OR4_154_Y, 
        OR4_238_Y, OR4_37_Y, OR4_32_Y, OR2_20_Y, OR4_187_Y, OR4_98_Y, 
        OR4_79_Y, OR4_68_Y, OR4_305_Y, OR4_233_Y, OR4_227_Y, OR4_93_Y, 
        OR4_21_Y, OR2_10_Y, OR4_246_Y, OR4_88_Y, OR4_142_Y, OR4_162_Y, 
        OR4_57_Y, OR4_317_Y, OR4_333_Y, OR4_31_Y, OR4_164_Y, OR2_37_Y, 
        OR4_342_Y, OR4_210_Y, OR4_23_Y, OR4_185_Y, OR4_286_Y, 
        OR4_359_Y, OR4_30_Y, OR4_300_Y, OR4_309_Y, OR2_12_Y, OR4_193_Y, 
        OR4_122_Y, OR4_95_Y, OR4_22_Y, OR4_341_Y, OR4_107_Y, OR4_253_Y, 
        OR4_38_Y, OR4_277_Y, OR2_32_Y, CFG3_6_Y, CFG3_0_Y, CFG3_8_Y, 
        CFG3_19_Y, CFG3_21_Y, CFG3_12_Y, CFG3_2_Y, CFG3_15_Y, CFG3_5_Y, 
        CFG3_17_Y, CFG3_9_Y, CFG3_22_Y, OR4_310_Y, OR4_264_Y, 
        OR4_105_Y, OR4_143_Y, OR4_198_Y, OR4_131_Y, OR4_65_Y, OR4_85_Y, 
        OR4_74_Y, OR2_27_Y, OR4_345_Y, OR4_330_Y, OR4_282_Y, OR4_124_Y, 
        OR4_42_Y, OR4_257_Y, OR4_332_Y, OR4_147_Y, OR4_172_Y, OR2_6_Y, 
        OR4_82_Y, OR4_251_Y, OR4_11_Y, OR4_55_Y, OR4_43_Y, OR4_158_Y, 
        OR4_90_Y, OR4_87_Y, OR4_69_Y, OR2_8_Y, OR4_27_Y, OR4_204_Y, 
        OR4_352_Y, OR4_242_Y, OR4_168_Y, OR4_18_Y, OR4_34_Y, OR4_218_Y, 
        OR4_64_Y, OR2_14_Y, OR4_328_Y, OR4_311_Y, OR4_320_Y, OR4_202_Y, 
        OR4_94_Y, OR4_146_Y, OR4_145_Y, OR4_207_Y, OR4_52_Y, OR2_29_Y, 
        OR4_294_Y, OR4_13_Y, OR4_171_Y, OR4_33_Y, OR4_266_Y, OR4_186_Y, 
        OR4_270_Y, OR4_73_Y, OR4_67_Y, OR2_4_Y, OR4_278_Y, OR4_66_Y, 
        OR4_121_Y, OR4_149_Y, OR4_35_Y, OR4_111_Y, OR4_39_Y, OR4_226_Y, 
        OR4_20_Y, OR2_31_Y, OR4_212_Y, OR4_130_Y, OR4_114_Y, OR4_106_Y, 
        OR4_336_Y, OR4_268_Y, OR4_258_Y, OR4_126_Y, OR4_53_Y, OR2_38_Y, 
        OR4_344_Y, OR4_295_Y, OR4_132_Y, OR4_173_Y, OR4_228_Y, 
        OR4_150_Y, OR4_102_Y, OR4_120_Y, OR4_108_Y, OR2_13_Y, OR4_0_Y, 
        OR4_346_Y, OR4_356_Y, OR4_237_Y, OR4_127_Y, OR4_178_Y, 
        OR4_177_Y, OR4_241_Y, OR4_92_Y, OR2_15_Y, CFG3_11_Y, CFG3_1_Y, 
        CFG3_16_Y, CFG3_23_Y, CFG3_18_Y, CFG3_14_Y, CFG3_7_Y, CFG3_3_Y, 
        CFG3_4_Y, CFG3_20_Y, CFG3_13_Y, CFG3_10_Y, OR4_58_Y, OR4_299_Y, 
        OR4_119_Y, OR4_271_Y, OR4_5_Y, OR4_80_Y, OR4_125_Y, OR4_17_Y, 
        OR4_25_Y, OR2_17_Y, VCC, GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    OR4 OR4_253 (.A(\R_DATA_TEMPR8[39] ), .B(\R_DATA_TEMPR9[39] ), .C(
        \R_DATA_TEMPR10[39] ), .D(\R_DATA_TEMPR11[39] ), .Y(OR4_253_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R29C2 (.BLK_EN(\BLKX0[29] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[29] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][2] ), .R_DATA({nc0, nc1, 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR29[28] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR29[26] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR29[24] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR29[22] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR29[20] }));
    OR4 OR4_181 (.A(OR4_284_Y), .B(OR2_26_Y), .C(\R_DATA_TEMPR22[24] ), 
        .D(\R_DATA_TEMPR23[24] ), .Y(OR4_181_Y));
    OR4 OR4_106 (.A(\R_DATA_TEMPR28[13] ), .B(\R_DATA_TEMPR29[13] ), 
        .C(\R_DATA_TEMPR30[13] ), .D(\R_DATA_TEMPR31[13] ), .Y(
        OR4_106_Y));
    OR4 OR4_83 (.A(OR4_201_Y), .B(OR4_267_Y), .C(OR4_265_Y), .D(
        OR4_323_Y), .Y(OR4_83_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[22]  (.A(CFG3_7_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[22] ));
    OR4 OR4_138 (.A(\R_DATA_TEMPR8[29] ), .B(\R_DATA_TEMPR9[29] ), .C(
        \R_DATA_TEMPR10[29] ), .D(\R_DATA_TEMPR11[29] ), .Y(OR4_138_Y));
    OR4 OR4_176 (.A(\R_DATA_TEMPR28[33] ), .B(\R_DATA_TEMPR29[33] ), 
        .C(\R_DATA_TEMPR30[33] ), .D(\R_DATA_TEMPR31[33] ), .Y(
        OR4_176_Y));
    OR4 OR4_308 (.A(OR4_249_Y), .B(OR4_327_Y), .C(OR4_8_Y), .D(
        OR4_273_Y), .Y(OR4_308_Y));
    OR4 OR4_317 (.A(\R_DATA_TEMPR4[36] ), .B(\R_DATA_TEMPR5[36] ), .C(
        \R_DATA_TEMPR6[36] ), .D(\R_DATA_TEMPR7[36] ), .Y(OR4_317_Y));
    OR4 OR4_110 (.A(\R_DATA_TEMPR0[3] ), .B(\R_DATA_TEMPR1[3] ), .C(
        \R_DATA_TEMPR2[3] ), .D(\R_DATA_TEMPR3[3] ), .Y(OR4_110_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_16 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_16_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R18C2 (.BLK_EN(\BLKX0[18] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][2] ), .R_DATA({nc2, nc3, 
        \R_DATA_TEMPR18[29] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR18[27] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR18[25] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR18[23] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR18[21] , \R_DATA_TEMPR18[20] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R7C3 (.BLK_EN(\BLKX0[7] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][3] ), .R_DATA({nc4, nc5, 
        \R_DATA_TEMPR7[39] , \R_DATA_TEMPR7[38] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR7[36] , \R_DATA_TEMPR7[35] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR7[33] , \R_DATA_TEMPR7[32] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR7[30] }));
    OR4 OR4_2 (.A(OR4_91_Y), .B(OR2_33_Y), .C(\R_DATA_TEMPR22[16] ), 
        .D(\R_DATA_TEMPR23[16] ), .Y(OR4_2_Y));
    OR4 OR4_329 (.A(OR4_281_Y), .B(OR2_30_Y), .C(\R_DATA_TEMPR22[37] ), 
        .D(\R_DATA_TEMPR23[37] ), .Y(OR4_329_Y));
    OR4 \OR4_R_DATA[29]  (.A(OR4_84_Y), .B(OR4_3_Y), .C(OR4_338_Y), .D(
        OR4_280_Y), .Y(R_DATA[29]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R4C2 (.BLK_EN(\BLKX0[4] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][2] ), .R_DATA({nc6, nc7, 
        \R_DATA_TEMPR4[29] , \R_DATA_TEMPR4[28] , \R_DATA_TEMPR4[27] , 
        \R_DATA_TEMPR4[26] , \R_DATA_TEMPR4[25] , \R_DATA_TEMPR4[24] , 
        \R_DATA_TEMPR4[23] , \R_DATA_TEMPR4[22] , \R_DATA_TEMPR4[21] , 
        \R_DATA_TEMPR4[20] }));
    OR4 OR4_48 (.A(\R_DATA_TEMPR28[26] ), .B(\R_DATA_TEMPR29[26] ), .C(
        \R_DATA_TEMPR30[26] ), .D(\R_DATA_TEMPR31[26] ), .Y(OR4_48_Y));
    OR4 OR4_109 (.A(\R_DATA_TEMPR0[17] ), .B(\R_DATA_TEMPR1[17] ), .C(
        \R_DATA_TEMPR2[17] ), .D(\R_DATA_TEMPR3[17] ), .Y(OR4_109_Y));
    OR2 OR2_33 (.A(\R_DATA_TEMPR20[16] ), .B(\R_DATA_TEMPR21[16] ), .Y(
        OR2_33_Y));
    OR2 OR2_15 (.A(\R_DATA_TEMPR20[11] ), .B(\R_DATA_TEMPR21[11] ), .Y(
        OR2_15_Y));
    OR4 OR4_241 (.A(\R_DATA_TEMPR12[11] ), .B(\R_DATA_TEMPR13[11] ), 
        .C(\R_DATA_TEMPR14[11] ), .D(\R_DATA_TEMPR15[11] ), .Y(
        OR4_241_Y));
    OR4 OR4_81 (.A(\R_DATA_TEMPR8[17] ), .B(\R_DATA_TEMPR9[17] ), .C(
        \R_DATA_TEMPR10[17] ), .D(\R_DATA_TEMPR11[17] ), .Y(OR4_81_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[29]  (.A(CFG3_14_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[29] ));
    OR4 OR4_118 (.A(OR4_182_Y), .B(OR2_3_Y), .C(\R_DATA_TEMPR22[9] ), 
        .D(\R_DATA_TEMPR23[9] ), .Y(OR4_118_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_206_Y), .B(OR4_325_Y), .C(OR4_224_Y), 
        .D(OR4_167_Y), .Y(R_DATA[7]));
    OR4 OR4_179 (.A(\R_DATA_TEMPR28[3] ), .B(\R_DATA_TEMPR29[3] ), .C(
        \R_DATA_TEMPR30[3] ), .D(\R_DATA_TEMPR31[3] ), .Y(OR4_179_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R26C1 (.BLK_EN(\BLKX0[26] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[26] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][1] ), .R_DATA({nc8, nc9, 
        \R_DATA_TEMPR26[19] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR26[17] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR26[15] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR26[13] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR26[11] , \R_DATA_TEMPR26[10] }));
    OR4 \OR4_R_DATA[4]  (.A(OR4_278_Y), .B(OR4_66_Y), .C(OR4_121_Y), 
        .D(OR4_149_Y), .Y(R_DATA[4]));
    OR4 OR4_135 (.A(OR4_307_Y), .B(OR4_199_Y), .C(OR4_217_Y), .D(
        OR4_289_Y), .Y(OR4_135_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[27]  (.A(CFG3_23_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[27] ));
    OR2 OR2_31 (.A(\R_DATA_TEMPR20[4] ), .B(\R_DATA_TEMPR21[4] ), .Y(
        OR2_31_Y));
    OR4 OR4_267 (.A(\R_DATA_TEMPR4[31] ), .B(\R_DATA_TEMPR5[31] ), .C(
        \R_DATA_TEMPR6[31] ), .D(\R_DATA_TEMPR7[31] ), .Y(OR4_267_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_9 (.A(BLK_EN), .B(R_ADDR[10]), .C(
        R_ADDR[9]), .Y(CFG3_9_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[4]  (.A(CFG3_18_Y), .B(CFG3_4_Y)
        , .Y(\BLKZ0[4] ));
    OR4 OR4_167 (.A(\R_DATA_TEMPR28[7] ), .B(\R_DATA_TEMPR29[7] ), .C(
        \R_DATA_TEMPR30[7] ), .D(\R_DATA_TEMPR31[7] ), .Y(OR4_167_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R6C3 (.BLK_EN(\BLKX0[6] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][3] ), .R_DATA({nc10, nc11, 
        \R_DATA_TEMPR6[39] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR6[37] , 
        \R_DATA_TEMPR6[36] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR6[34] , 
        \R_DATA_TEMPR6[33] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR6[31] , 
        \R_DATA_TEMPR6[30] }));
    OR4 OR4_186 (.A(\R_DATA_TEMPR4[10] ), .B(\R_DATA_TEMPR5[10] ), .C(
        \R_DATA_TEMPR6[10] ), .D(\R_DATA_TEMPR7[10] ), .Y(OR4_186_Y));
    OR4 OR4_341 (.A(\R_DATA_TEMPR0[39] ), .B(\R_DATA_TEMPR1[39] ), .C(
        \R_DATA_TEMPR2[39] ), .D(\R_DATA_TEMPR3[39] ), .Y(OR4_341_Y));
    OR4 OR4_235 (.A(\R_DATA_TEMPR16[8] ), .B(\R_DATA_TEMPR17[8] ), .C(
        \R_DATA_TEMPR18[8] ), .D(\R_DATA_TEMPR19[8] ), .Y(OR4_235_Y));
    OR2 OR2_29 (.A(\R_DATA_TEMPR20[21] ), .B(\R_DATA_TEMPR21[21] ), .Y(
        OR2_29_Y));
    OR4 OR4_264 (.A(OR4_74_Y), .B(OR2_27_Y), .C(\R_DATA_TEMPR22[28] ), 
        .D(\R_DATA_TEMPR23[28] ), .Y(OR4_264_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R4C0 (.BLK_EN(\BLKX0[4] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][0] ), .R_DATA({nc12, nc13, 
        \R_DATA_TEMPR4[9] , \R_DATA_TEMPR4[8] , \R_DATA_TEMPR4[7] , 
        \R_DATA_TEMPR4[6] , \R_DATA_TEMPR4[5] , \R_DATA_TEMPR4[4] , 
        \R_DATA_TEMPR4[3] , \R_DATA_TEMPR4[2] , \R_DATA_TEMPR4[1] , 
        \R_DATA_TEMPR4[0] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R23C0 (.BLK_EN(\BLKX0[23] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[23] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][0] ), .R_DATA({nc14, nc15, 
        \R_DATA_TEMPR23[9] , \R_DATA_TEMPR23[8] , \R_DATA_TEMPR23[7] , 
        \R_DATA_TEMPR23[6] , \R_DATA_TEMPR23[5] , \R_DATA_TEMPR23[4] , 
        \R_DATA_TEMPR23[3] , \R_DATA_TEMPR23[2] , \R_DATA_TEMPR23[1] , 
        \R_DATA_TEMPR23[0] }));
    OR4 OR4_293 (.A(\R_DATA_TEMPR28[0] ), .B(\R_DATA_TEMPR29[0] ), .C(
        \R_DATA_TEMPR30[0] ), .D(\R_DATA_TEMPR31[0] ), .Y(OR4_293_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[15]  (.A(CFG3_15_Y), .B(
        CFG3_17_Y), .Y(\BLKX0[15] ));
    OR4 OR4_115 (.A(\R_DATA_TEMPR12[25] ), .B(\R_DATA_TEMPR13[25] ), 
        .C(\R_DATA_TEMPR14[25] ), .D(\R_DATA_TEMPR15[25] ), .Y(
        OR4_115_Y));
    OR4 OR4_66 (.A(OR4_20_Y), .B(OR2_31_Y), .C(\R_DATA_TEMPR22[4] ), 
        .D(\R_DATA_TEMPR23[4] ), .Y(OR4_66_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[10]  (.A(CFG3_16_Y), .B(
        CFG3_20_Y), .Y(\BLKZ0[10] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[8]  (.A(CFG3_6_Y), .B(CFG3_17_Y)
        , .Y(\BLKX0[8] ));
    OR4 OR4_238 (.A(\R_DATA_TEMPR8[20] ), .B(\R_DATA_TEMPR9[20] ), .C(
        \R_DATA_TEMPR10[20] ), .D(\R_DATA_TEMPR11[20] ), .Y(OR4_238_Y));
    OR2 OR2_8 (.A(\R_DATA_TEMPR20[6] ), .B(\R_DATA_TEMPR21[6] ), .Y(
        OR2_8_Y));
    OR4 OR4_189 (.A(\R_DATA_TEMPR16[19] ), .B(\R_DATA_TEMPR17[19] ), 
        .C(\R_DATA_TEMPR18[19] ), .D(\R_DATA_TEMPR19[19] ), .Y(
        OR4_189_Y));
    OR4 OR4_0 (.A(OR4_127_Y), .B(OR4_178_Y), .C(OR4_177_Y), .D(
        OR4_241_Y), .Y(OR4_0_Y));
    OR4 OR4_207 (.A(\R_DATA_TEMPR12[21] ), .B(\R_DATA_TEMPR13[21] ), 
        .C(\R_DATA_TEMPR14[21] ), .D(\R_DATA_TEMPR15[21] ), .Y(
        OR4_207_Y));
    OR4 OR4_215 (.A(\R_DATA_TEMPR12[7] ), .B(\R_DATA_TEMPR13[7] ), .C(
        \R_DATA_TEMPR14[7] ), .D(\R_DATA_TEMPR15[7] ), .Y(OR4_215_Y));
    OR4 OR4_107 (.A(\R_DATA_TEMPR4[39] ), .B(\R_DATA_TEMPR5[39] ), .C(
        \R_DATA_TEMPR6[39] ), .D(\R_DATA_TEMPR7[39] ), .Y(OR4_107_Y));
    OR4 OR4_277 (.A(\R_DATA_TEMPR16[39] ), .B(\R_DATA_TEMPR17[39] ), 
        .C(\R_DATA_TEMPR18[39] ), .D(\R_DATA_TEMPR19[39] ), .Y(
        OR4_277_Y));
    OR4 OR4_95 (.A(\R_DATA_TEMPR24[39] ), .B(\R_DATA_TEMPR25[39] ), .C(
        \R_DATA_TEMPR26[39] ), .D(\R_DATA_TEMPR27[39] ), .Y(OR4_95_Y));
    OR2 OR2_22 (.A(\R_DATA_TEMPR20[25] ), .B(\R_DATA_TEMPR21[25] ), .Y(
        OR2_22_Y));
    OR4 OR4_177 (.A(\R_DATA_TEMPR8[11] ), .B(\R_DATA_TEMPR9[11] ), .C(
        \R_DATA_TEMPR10[11] ), .D(\R_DATA_TEMPR11[11] ), .Y(OR4_177_Y));
    OR4 \OR4_R_DATA[34]  (.A(OR4_58_Y), .B(OR4_299_Y), .C(OR4_119_Y), 
        .D(OR4_271_Y), .Y(R_DATA[34]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R5C1 (.BLK_EN(\BLKX0[5] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][1] ), .R_DATA({nc16, nc17, 
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR5[18] , \R_DATA_TEMPR5[17] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR5[15] , \R_DATA_TEMPR5[14] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR5[12] , \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR5[10] }));
    OR4 OR4_349 (.A(\R_DATA_TEMPR16[15] ), .B(\R_DATA_TEMPR17[15] ), 
        .C(\R_DATA_TEMPR18[15] ), .D(\R_DATA_TEMPR19[15] ), .Y(
        OR4_349_Y));
    OR4 OR4_223 (.A(\R_DATA_TEMPR0[29] ), .B(\R_DATA_TEMPR1[29] ), .C(
        \R_DATA_TEMPR2[29] ), .D(\R_DATA_TEMPR3[29] ), .Y(OR4_223_Y));
    OR4 OR4_354 (.A(\R_DATA_TEMPR0[30] ), .B(\R_DATA_TEMPR1[30] ), .C(
        \R_DATA_TEMPR2[30] ), .D(\R_DATA_TEMPR3[30] ), .Y(OR4_354_Y));
    OR4 OR4_204 (.A(OR4_64_Y), .B(OR2_14_Y), .C(\R_DATA_TEMPR22[35] ), 
        .D(\R_DATA_TEMPR23[35] ), .Y(OR4_204_Y));
    OR2 OR2_19 (.A(\R_DATA_TEMPR20[31] ), .B(\R_DATA_TEMPR21[31] ), .Y(
        OR2_19_Y));
    OR4 OR4_151 (.A(\R_DATA_TEMPR24[3] ), .B(\R_DATA_TEMPR25[3] ), .C(
        \R_DATA_TEMPR26[3] ), .D(\R_DATA_TEMPR27[3] ), .Y(OR4_151_Y));
    OR4 OR4_274 (.A(\R_DATA_TEMPR28[2] ), .B(\R_DATA_TEMPR29[2] ), .C(
        \R_DATA_TEMPR30[2] ), .D(\R_DATA_TEMPR31[2] ), .Y(OR4_274_Y));
    OR4 OR4_218 (.A(\R_DATA_TEMPR12[35] ), .B(\R_DATA_TEMPR13[35] ), 
        .C(\R_DATA_TEMPR14[35] ), .D(\R_DATA_TEMPR15[35] ), .Y(
        OR4_218_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_225_Y), .B(OR4_213_Y), .C(OR4_163_Y), 
        .D(OR4_7_Y), .Y(R_DATA[22]));
    OR4 OR4_60 (.A(OR4_314_Y), .B(OR4_239_Y), .C(OR4_175_Y), .D(
        OR4_194_Y), .Y(OR4_60_Y));
    OR4 OR4_67 (.A(\R_DATA_TEMPR16[10] ), .B(\R_DATA_TEMPR17[10] ), .C(
        \R_DATA_TEMPR18[10] ), .D(\R_DATA_TEMPR19[10] ), .Y(OR4_67_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R23C3 (.BLK_EN(\BLKX0[23] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[23] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][3] ), .R_DATA({nc18, nc19, 
        \R_DATA_TEMPR23[39] , \R_DATA_TEMPR23[38] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR23[36] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR23[34] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR23[32] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR23[30] }));
    OR4 OR4_305 (.A(\R_DATA_TEMPR0[23] ), .B(\R_DATA_TEMPR1[23] ), .C(
        \R_DATA_TEMPR2[23] ), .D(\R_DATA_TEMPR3[23] ), .Y(OR4_305_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[0]  (.A(CFG3_6_Y), .B(CFG3_5_Y), 
        .Y(\BLKX0[0] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[13]  (.A(CFG3_14_Y), .B(
        CFG3_20_Y), .Y(\BLKZ0[13] ));
    OR4 OR4_232 (.A(\R_DATA_TEMPR0[20] ), .B(\R_DATA_TEMPR1[20] ), .C(
        \R_DATA_TEMPR2[20] ), .D(\R_DATA_TEMPR3[20] ), .Y(OR4_232_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_6 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_6_Y));
    OR4 \OR4_R_DATA[15]  (.A(OR4_312_Y), .B(OR4_129_Y), .C(OR4_263_Y), 
        .D(OR4_156_Y), .Y(R_DATA[15]));
    OR4 OR4_45 (.A(\R_DATA_TEMPR8[27] ), .B(\R_DATA_TEMPR9[27] ), .C(
        \R_DATA_TEMPR10[27] ), .D(\R_DATA_TEMPR11[27] ), .Y(OR4_45_Y));
    OR4 OR4_160 (.A(OR4_340_Y), .B(OR4_229_Y), .C(OR4_248_Y), .D(
        OR4_318_Y), .Y(OR4_160_Y));
    OR2 OR2_12 (.A(\R_DATA_TEMPR20[14] ), .B(\R_DATA_TEMPR21[14] ), .Y(
        OR2_12_Y));
    OR4 \OR4_R_DATA[23]  (.A(OR4_187_Y), .B(OR4_98_Y), .C(OR4_79_Y), 
        .D(OR4_68_Y), .Y(R_DATA[23]));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[26]  (.A(CFG3_8_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[26] ));
    OR4 OR4_330 (.A(OR4_172_Y), .B(OR2_6_Y), .C(\R_DATA_TEMPR22[32] ), 
        .D(\R_DATA_TEMPR23[32] ), .Y(OR4_330_Y));
    OR4 OR4_287 (.A(\R_DATA_TEMPR0[0] ), .B(\R_DATA_TEMPR1[0] ), .C(
        \R_DATA_TEMPR2[0] ), .D(\R_DATA_TEMPR3[0] ), .Y(OR4_287_Y));
    OR4 OR4_86 (.A(\R_DATA_TEMPR28[16] ), .B(\R_DATA_TEMPR29[16] ), .C(
        \R_DATA_TEMPR30[16] ), .D(\R_DATA_TEMPR31[16] ), .Y(OR4_86_Y));
    OR4 OR4_33 (.A(\R_DATA_TEMPR28[10] ), .B(\R_DATA_TEMPR29[10] ), .C(
        \R_DATA_TEMPR30[10] ), .D(\R_DATA_TEMPR31[10] ), .Y(OR4_33_Y));
    OR4 OR4_168 (.A(\R_DATA_TEMPR0[35] ), .B(\R_DATA_TEMPR1[35] ), .C(
        \R_DATA_TEMPR2[35] ), .D(\R_DATA_TEMPR3[35] ), .Y(OR4_168_Y));
    OR4 OR4_187 (.A(OR4_305_Y), .B(OR4_233_Y), .C(OR4_227_Y), .D(
        OR4_93_Y), .Y(OR4_187_Y));
    OR4 OR4_212 (.A(OR4_336_Y), .B(OR4_268_Y), .C(OR4_258_Y), .D(
        OR4_126_Y), .Y(OR4_212_Y));
    OR4 OR4_353 (.A(\R_DATA_TEMPR12[0] ), .B(\R_DATA_TEMPR13[0] ), .C(
        \R_DATA_TEMPR14[0] ), .D(\R_DATA_TEMPR15[0] ), .Y(OR4_353_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R15C0 (.BLK_EN(\BLKX0[15] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][0] ), .R_DATA({nc20, nc21, 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR15[0] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[6]  (.A(CFG3_2_Y), .B(CFG3_5_Y), 
        .Y(\BLKX0[6] ));
    OR4 OR4_284 (.A(\R_DATA_TEMPR16[24] ), .B(\R_DATA_TEMPR17[24] ), 
        .C(\R_DATA_TEMPR18[24] ), .D(\R_DATA_TEMPR19[24] ), .Y(
        OR4_284_Y));
    OR4 OR4_310 (.A(OR4_198_Y), .B(OR4_131_Y), .C(OR4_65_Y), .D(
        OR4_85_Y), .Y(OR4_310_Y));
    OR4 OR4_5 (.A(\R_DATA_TEMPR0[34] ), .B(\R_DATA_TEMPR1[34] ), .C(
        \R_DATA_TEMPR2[34] ), .D(\R_DATA_TEMPR3[34] ), .Y(OR4_5_Y));
    OR4 OR4_307 (.A(\R_DATA_TEMPR0[26] ), .B(\R_DATA_TEMPR1[26] ), .C(
        \R_DATA_TEMPR2[26] ), .D(\R_DATA_TEMPR3[26] ), .Y(OR4_307_Y));
    OR4 OR4_100 (.A(\R_DATA_TEMPR16[12] ), .B(\R_DATA_TEMPR17[12] ), 
        .C(\R_DATA_TEMPR18[12] ), .D(\R_DATA_TEMPR19[12] ), .Y(
        OR4_100_Y));
    OR4 OR4_99 (.A(\R_DATA_TEMPR28[37] ), .B(\R_DATA_TEMPR29[37] ), .C(
        \R_DATA_TEMPR30[37] ), .D(\R_DATA_TEMPR31[37] ), .Y(OR4_99_Y));
    OR4 OR4_156 (.A(\R_DATA_TEMPR28[15] ), .B(\R_DATA_TEMPR29[15] ), 
        .C(\R_DATA_TEMPR30[15] ), .D(\R_DATA_TEMPR31[15] ), .Y(
        OR4_156_Y));
    OR2 OR2_36 (.A(\R_DATA_TEMPR20[27] ), .B(\R_DATA_TEMPR21[27] ), .Y(
        OR2_36_Y));
    OR4 OR4_68 (.A(\R_DATA_TEMPR28[23] ), .B(\R_DATA_TEMPR29[23] ), .C(
        \R_DATA_TEMPR30[23] ), .D(\R_DATA_TEMPR31[23] ), .Y(OR4_68_Y));
    OR2 OR2_24 (.A(\R_DATA_TEMPR20[17] ), .B(\R_DATA_TEMPR21[17] ), .Y(
        OR2_24_Y));
    OR4 OR4_170 (.A(OR4_240_Y), .B(OR2_23_Y), .C(\R_DATA_TEMPR22[2] ), 
        .D(\R_DATA_TEMPR23[2] ), .Y(OR4_170_Y));
    OR4 OR4_31 (.A(\R_DATA_TEMPR12[36] ), .B(\R_DATA_TEMPR13[36] ), .C(
        \R_DATA_TEMPR14[36] ), .D(\R_DATA_TEMPR15[36] ), .Y(OR4_31_Y));
    OR4 \OR4_R_DATA[31]  (.A(OR4_83_Y), .B(OR4_61_Y), .C(OR4_70_Y), .D(
        OR4_321_Y), .Y(R_DATA[31]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R16C2 (.BLK_EN(\BLKX0[16] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][2] ), .R_DATA({nc22, nc23, 
        \R_DATA_TEMPR16[29] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR16[27] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR16[25] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR16[23] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR16[21] , \R_DATA_TEMPR16[20] }));
    OR4 OR4_243 (.A(\R_DATA_TEMPR24[2] ), .B(\R_DATA_TEMPR25[2] ), .C(
        \R_DATA_TEMPR26[2] ), .D(\R_DATA_TEMPR27[2] ), .Y(OR4_243_Y));
    OR4 OR4_358 (.A(\R_DATA_TEMPR8[30] ), .B(\R_DATA_TEMPR9[30] ), .C(
        \R_DATA_TEMPR10[30] ), .D(\R_DATA_TEMPR11[30] ), .Y(OR4_358_Y));
    OR4 OR4_80 (.A(\R_DATA_TEMPR4[34] ), .B(\R_DATA_TEMPR5[34] ), .C(
        \R_DATA_TEMPR6[34] ), .D(\R_DATA_TEMPR7[34] ), .Y(OR4_80_Y));
    OR4 OR4_108 (.A(\R_DATA_TEMPR16[18] ), .B(\R_DATA_TEMPR17[18] ), 
        .C(\R_DATA_TEMPR18[18] ), .D(\R_DATA_TEMPR19[18] ), .Y(
        OR4_108_Y));
    OR4 OR4_191 (.A(\R_DATA_TEMPR24[33] ), .B(\R_DATA_TEMPR25[33] ), 
        .C(\R_DATA_TEMPR26[33] ), .D(\R_DATA_TEMPR27[33] ), .Y(
        OR4_191_Y));
    OR4 OR4_1 (.A(\R_DATA_TEMPR24[24] ), .B(\R_DATA_TEMPR25[24] ), .C(
        \R_DATA_TEMPR26[24] ), .D(\R_DATA_TEMPR27[24] ), .Y(OR4_1_Y));
    OR4 OR4_87 (.A(\R_DATA_TEMPR12[6] ), .B(\R_DATA_TEMPR13[6] ), .C(
        \R_DATA_TEMPR14[6] ), .D(\R_DATA_TEMPR15[6] ), .Y(OR4_87_Y));
    OR4 \OR4_R_DATA[30]  (.A(OR4_14_Y), .B(OR4_103_Y), .C(OR4_259_Y), 
        .D(OR4_128_Y), .Y(R_DATA[30]));
    OR4 OR4_178 (.A(\R_DATA_TEMPR4[11] ), .B(\R_DATA_TEMPR5[11] ), .C(
        \R_DATA_TEMPR6[11] ), .D(\R_DATA_TEMPR7[11] ), .Y(OR4_178_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R26C0 (.BLK_EN(\BLKX0[26] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[26] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][0] ), .R_DATA({nc24, nc25, 
        \R_DATA_TEMPR26[9] , \R_DATA_TEMPR26[8] , \R_DATA_TEMPR26[7] , 
        \R_DATA_TEMPR26[6] , \R_DATA_TEMPR26[5] , \R_DATA_TEMPR26[4] , 
        \R_DATA_TEMPR26[3] , \R_DATA_TEMPR26[2] , \R_DATA_TEMPR26[1] , 
        \R_DATA_TEMPR26[0] }));
    OR4 OR4_159 (.A(\R_DATA_TEMPR8[37] ), .B(\R_DATA_TEMPR9[37] ), .C(
        \R_DATA_TEMPR10[37] ), .D(\R_DATA_TEMPR11[37] ), .Y(OR4_159_Y));
    OR4 OR4_165 (.A(\R_DATA_TEMPR16[31] ), .B(\R_DATA_TEMPR17[31] ), 
        .C(\R_DATA_TEMPR18[31] ), .D(\R_DATA_TEMPR19[31] ), .Y(
        OR4_165_Y));
    OR4 OR4_133 (.A(\R_DATA_TEMPR28[25] ), .B(\R_DATA_TEMPR29[25] ), 
        .C(\R_DATA_TEMPR30[25] ), .D(\R_DATA_TEMPR31[25] ), .Y(
        OR4_133_Y));
    OR4 OR4_92 (.A(\R_DATA_TEMPR16[11] ), .B(\R_DATA_TEMPR17[11] ), .C(
        \R_DATA_TEMPR18[11] ), .D(\R_DATA_TEMPR19[11] ), .Y(OR4_92_Y));
    OR4 \OR4_R_DATA[36]  (.A(OR4_246_Y), .B(OR4_88_Y), .C(OR4_142_Y), 
        .D(OR4_162_Y), .Y(R_DATA[36]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R4C3 (.BLK_EN(\BLKX0[4] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][3] ), .R_DATA({nc26, nc27, 
        \R_DATA_TEMPR4[39] , \R_DATA_TEMPR4[38] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR4[36] , \R_DATA_TEMPR4[35] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR4[33] , \R_DATA_TEMPR4[32] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR4[30] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[11]  (.A(CFG3_23_Y), .B(
        CFG3_20_Y), .Y(\BLKZ0[11] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[16]  (.A(CFG3_11_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[16] ));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R18C1 (.BLK_EN(\BLKX0[18] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][1] ), .R_DATA({nc28, nc29, 
        \R_DATA_TEMPR18[19] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR18[17] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR18[15] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR18[13] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR18[11] , \R_DATA_TEMPR18[10] }));
    OR2 OR2_30 (.A(\R_DATA_TEMPR20[37] ), .B(\R_DATA_TEMPR21[37] ), .Y(
        OR2_30_Y));
    OR4 OR4_324 (.A(\R_DATA_TEMPR0[12] ), .B(\R_DATA_TEMPR1[12] ), .C(
        \R_DATA_TEMPR2[12] ), .D(\R_DATA_TEMPR3[12] ), .Y(OR4_324_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R28C0 (.BLK_EN(\BLKX0[28] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[28] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][0] ), .R_DATA({nc30, nc31, 
        \R_DATA_TEMPR28[9] , \R_DATA_TEMPR28[8] , \R_DATA_TEMPR28[7] , 
        \R_DATA_TEMPR28[6] , \R_DATA_TEMPR28[5] , \R_DATA_TEMPR28[4] , 
        \R_DATA_TEMPR28[3] , \R_DATA_TEMPR28[2] , \R_DATA_TEMPR28[1] , 
        \R_DATA_TEMPR28[0] }));
    OR4 OR4_265 (.A(\R_DATA_TEMPR8[31] ), .B(\R_DATA_TEMPR9[31] ), .C(
        \R_DATA_TEMPR10[31] ), .D(\R_DATA_TEMPR11[31] ), .Y(OR4_265_Y));
    OR4 OR4_49 (.A(\R_DATA_TEMPR16[26] ), .B(\R_DATA_TEMPR17[26] ), .C(
        \R_DATA_TEMPR18[26] ), .D(\R_DATA_TEMPR19[26] ), .Y(OR4_49_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R4C1 (.BLK_EN(\BLKX0[4] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][1] ), .R_DATA({nc32, nc33, 
        \R_DATA_TEMPR4[19] , \R_DATA_TEMPR4[18] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR4[16] , \R_DATA_TEMPR4[15] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR4[13] , \R_DATA_TEMPR4[12] , \R_DATA_TEMPR4[11] , 
        \R_DATA_TEMPR4[10] }));
    OR2 OR2_14 (.A(\R_DATA_TEMPR20[35] ), .B(\R_DATA_TEMPR21[35] ), .Y(
        OR2_14_Y));
    OR2 OR2_37 (.A(\R_DATA_TEMPR20[36] ), .B(\R_DATA_TEMPR21[36] ), .Y(
        OR2_37_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R19C2 (.BLK_EN(\BLKX0[19] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][2] ), .R_DATA({nc34, nc35, 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR19[28] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR19[26] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR19[24] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR19[22] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR19[20] }));
    OR4 OR4_121 (.A(\R_DATA_TEMPR24[4] ), .B(\R_DATA_TEMPR25[4] ), .C(
        \R_DATA_TEMPR26[4] ), .D(\R_DATA_TEMPR27[4] ), .Y(OR4_121_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R3C2 (.BLK_EN(\BLKX0[3] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][2] ), .R_DATA({nc36, nc37, 
        \R_DATA_TEMPR3[29] , \R_DATA_TEMPR3[28] , \R_DATA_TEMPR3[27] , 
        \R_DATA_TEMPR3[26] , \R_DATA_TEMPR3[25] , \R_DATA_TEMPR3[24] , 
        \R_DATA_TEMPR3[23] , \R_DATA_TEMPR3[22] , \R_DATA_TEMPR3[21] , 
        \R_DATA_TEMPR3[20] }));
    OR4 \OR4_R_DATA[18]  (.A(OR4_344_Y), .B(OR4_295_Y), .C(OR4_132_Y), 
        .D(OR4_173_Y), .Y(R_DATA[18]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R7C0 (.BLK_EN(\BLKX0[7] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][0] ), .R_DATA({nc38, nc39, 
        \R_DATA_TEMPR7[9] , \R_DATA_TEMPR7[8] , \R_DATA_TEMPR7[7] , 
        \R_DATA_TEMPR7[6] , \R_DATA_TEMPR7[5] , \R_DATA_TEMPR7[4] , 
        \R_DATA_TEMPR7[3] , \R_DATA_TEMPR7[2] , \R_DATA_TEMPR7[1] , 
        \R_DATA_TEMPR7[0] }));
    OR4 OR4_113 (.A(\R_DATA_TEMPR4[2] ), .B(\R_DATA_TEMPR5[2] ), .C(
        \R_DATA_TEMPR6[2] ), .D(\R_DATA_TEMPR7[2] ), .Y(OR4_113_Y));
    OR4 OR4_132 (.A(\R_DATA_TEMPR24[18] ), .B(\R_DATA_TEMPR25[18] ), 
        .C(\R_DATA_TEMPR26[18] ), .D(\R_DATA_TEMPR27[18] ), .Y(
        OR4_132_Y));
    OR4 OR4_7 (.A(\R_DATA_TEMPR28[22] ), .B(\R_DATA_TEMPR29[22] ), .C(
        \R_DATA_TEMPR30[22] ), .D(\R_DATA_TEMPR31[22] ), .Y(OR4_7_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[9]  (.A(CFG3_0_Y), .B(CFG3_17_Y)
        , .Y(\BLKX0[9] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[12]  (.A(CFG3_21_Y), .B(
        CFG3_17_Y), .Y(\BLKX0[12] ));
    OR4 OR4_268 (.A(\R_DATA_TEMPR4[13] ), .B(\R_DATA_TEMPR5[13] ), .C(
        \R_DATA_TEMPR6[13] ), .D(\R_DATA_TEMPR7[13] ), .Y(OR4_268_Y));
    OR4 OR4_180 (.A(OR4_139_Y), .B(OR2_9_Y), .C(\R_DATA_TEMPR22[3] ), 
        .D(\R_DATA_TEMPR23[3] ), .Y(OR4_180_Y));
    OR4 OR4_105 (.A(\R_DATA_TEMPR24[28] ), .B(\R_DATA_TEMPR25[28] ), 
        .C(\R_DATA_TEMPR26[28] ), .D(\R_DATA_TEMPR27[28] ), .Y(
        OR4_105_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[27]  (.A(CFG3_19_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[27] ));
    OR4 OR4_175 (.A(\R_DATA_TEMPR8[38] ), .B(\R_DATA_TEMPR9[38] ), .C(
        \R_DATA_TEMPR10[38] ), .D(\R_DATA_TEMPR11[38] ), .Y(OR4_175_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_15 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_15_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[1]  (.A(CFG3_1_Y), .B(CFG3_4_Y), 
        .Y(\BLKZ0[1] ));
    OR4 OR4_239 (.A(\R_DATA_TEMPR4[38] ), .B(\R_DATA_TEMPR5[38] ), .C(
        \R_DATA_TEMPR6[38] ), .D(\R_DATA_TEMPR7[38] ), .Y(OR4_239_Y));
    OR4 OR4_42 (.A(\R_DATA_TEMPR0[32] ), .B(\R_DATA_TEMPR1[32] ), .C(
        \R_DATA_TEMPR2[32] ), .D(\R_DATA_TEMPR3[32] ), .Y(OR4_42_Y));
    OR4 OR4_88 (.A(OR4_164_Y), .B(OR2_37_Y), .C(\R_DATA_TEMPR22[36] ), 
        .D(\R_DATA_TEMPR23[36] ), .Y(OR4_88_Y));
    OR4 OR4_205 (.A(OR4_137_Y), .B(OR2_1_Y), .C(\R_DATA_TEMPR22[33] ), 
        .D(\R_DATA_TEMPR23[33] ), .Y(OR4_205_Y));
    OR4 OR4_188 (.A(\R_DATA_TEMPR28[1] ), .B(\R_DATA_TEMPR29[1] ), .C(
        \R_DATA_TEMPR30[1] ), .D(\R_DATA_TEMPR31[1] ), .Y(OR4_188_Y));
    OR4 OR4_196 (.A(\R_DATA_TEMPR24[12] ), .B(\R_DATA_TEMPR25[12] ), 
        .C(\R_DATA_TEMPR26[12] ), .D(\R_DATA_TEMPR27[12] ), .Y(
        OR4_196_Y));
    OR4 OR4_112 (.A(\R_DATA_TEMPR12[5] ), .B(\R_DATA_TEMPR13[5] ), .C(
        \R_DATA_TEMPR14[5] ), .D(\R_DATA_TEMPR15[5] ), .Y(OR4_112_Y));
    OR4 OR4_275 (.A(\R_DATA_TEMPR4[25] ), .B(\R_DATA_TEMPR5[25] ), .C(
        \R_DATA_TEMPR6[25] ), .D(\R_DATA_TEMPR7[25] ), .Y(OR4_275_Y));
    OR4 \OR4_R_DATA[37]  (.A(OR4_153_Y), .B(OR4_329_Y), .C(OR4_56_Y), 
        .D(OR4_99_Y), .Y(R_DATA[37]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R16C1 (.BLK_EN(\BLKX0[16] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][1] ), .R_DATA({nc40, nc41, 
        \R_DATA_TEMPR16[19] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR16[17] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR16[15] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR16[13] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR16[11] , \R_DATA_TEMPR16[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R0C2 (.BLK_EN(\BLKX0[0] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][2] ), .R_DATA({nc42, nc43, 
        \R_DATA_TEMPR0[29] , \R_DATA_TEMPR0[28] , \R_DATA_TEMPR0[27] , 
        \R_DATA_TEMPR0[26] , \R_DATA_TEMPR0[25] , \R_DATA_TEMPR0[24] , 
        \R_DATA_TEMPR0[23] , \R_DATA_TEMPR0[22] , \R_DATA_TEMPR0[21] , 
        \R_DATA_TEMPR0[20] }));
    OR4 OR4_257 (.A(\R_DATA_TEMPR4[32] ), .B(\R_DATA_TEMPR5[32] ), .C(
        \R_DATA_TEMPR6[32] ), .D(\R_DATA_TEMPR7[32] ), .Y(OR4_257_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R27C3 (.BLK_EN(\BLKX0[27] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[27] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][3] ), .R_DATA({nc44, nc45, 
        \R_DATA_TEMPR27[39] , \R_DATA_TEMPR27[38] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR27[36] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR27[34] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR27[32] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR27[30] }));
    OR4 OR4_157 (.A(\R_DATA_TEMPR0[5] ), .B(\R_DATA_TEMPR1[5] ), .C(
        \R_DATA_TEMPR2[5] ), .D(\R_DATA_TEMPR3[5] ), .Y(OR4_157_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_7 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_7_Y));
    OR4 OR4_208 (.A(\R_DATA_TEMPR24[38] ), .B(\R_DATA_TEMPR25[38] ), 
        .C(\R_DATA_TEMPR26[38] ), .D(\R_DATA_TEMPR27[38] ), .Y(
        OR4_208_Y));
    OR4 OR4_219 (.A(\R_DATA_TEMPR12[27] ), .B(\R_DATA_TEMPR13[27] ), 
        .C(\R_DATA_TEMPR14[27] ), .D(\R_DATA_TEMPR15[27] ), .Y(
        OR4_219_Y));
    OR4 OR4_323 (.A(\R_DATA_TEMPR12[31] ), .B(\R_DATA_TEMPR13[31] ), 
        .C(\R_DATA_TEMPR14[31] ), .D(\R_DATA_TEMPR15[31] ), .Y(
        OR4_323_Y));
    OR4 \OR4_R_DATA[19]  (.A(OR4_117_Y), .B(OR4_26_Y), .C(OR4_9_Y), .D(
        OR4_304_Y), .Y(R_DATA[19]));
    OR2 OR2_38 (.A(\R_DATA_TEMPR20[13] ), .B(\R_DATA_TEMPR21[13] ), .Y(
        OR2_38_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R29C0 (.BLK_EN(\BLKX0[29] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[29] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][0] ), .R_DATA({nc46, nc47, 
        \R_DATA_TEMPR29[9] , \R_DATA_TEMPR29[8] , \R_DATA_TEMPR29[7] , 
        \R_DATA_TEMPR29[6] , \R_DATA_TEMPR29[5] , \R_DATA_TEMPR29[4] , 
        \R_DATA_TEMPR29[3] , \R_DATA_TEMPR29[2] , \R_DATA_TEMPR29[1] , 
        \R_DATA_TEMPR29[0] }));
    OR4 OR4_278 (.A(OR4_35_Y), .B(OR4_111_Y), .C(OR4_39_Y), .D(
        OR4_226_Y), .Y(OR4_278_Y));
    OR4 OR4_23 (.A(\R_DATA_TEMPR24[14] ), .B(\R_DATA_TEMPR25[14] ), .C(
        \R_DATA_TEMPR26[14] ), .D(\R_DATA_TEMPR27[14] ), .Y(OR4_23_Y));
    OR4 OR4_199 (.A(\R_DATA_TEMPR4[26] ), .B(\R_DATA_TEMPR5[26] ), .C(
        \R_DATA_TEMPR6[26] ), .D(\R_DATA_TEMPR7[26] ), .Y(OR4_199_Y));
    OR4 OR4_254 (.A(\R_DATA_TEMPR0[19] ), .B(\R_DATA_TEMPR1[19] ), .C(
        \R_DATA_TEMPR2[19] ), .D(\R_DATA_TEMPR3[19] ), .Y(OR4_254_Y));
    OR4 OR4_262 (.A(OR4_232_Y), .B(OR4_154_Y), .C(OR4_238_Y), .D(
        OR4_37_Y), .Y(OR4_262_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R29C3 (.BLK_EN(\BLKX0[29] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[29] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][3] ), .R_DATA({nc48, nc49, 
        \R_DATA_TEMPR29[39] , \R_DATA_TEMPR29[38] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR29[36] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR29[34] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR29[32] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR29[30] }));
    OR4 OR4_126 (.A(\R_DATA_TEMPR12[13] ), .B(\R_DATA_TEMPR13[13] ), 
        .C(\R_DATA_TEMPR14[13] ), .D(\R_DATA_TEMPR15[13] ), .Y(
        OR4_126_Y));
    OR4 OR4_94 (.A(\R_DATA_TEMPR0[21] ), .B(\R_DATA_TEMPR1[21] ), .C(
        \R_DATA_TEMPR2[21] ), .D(\R_DATA_TEMPR3[21] ), .Y(OR4_94_Y));
    OR4 OR4_65 (.A(\R_DATA_TEMPR8[28] ), .B(\R_DATA_TEMPR9[28] ), .C(
        \R_DATA_TEMPR10[28] ), .D(\R_DATA_TEMPR11[28] ), .Y(OR4_65_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R1C2 (.BLK_EN(\BLKX0[1] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][2] ), .R_DATA({nc50, nc51, 
        \R_DATA_TEMPR1[29] , \R_DATA_TEMPR1[28] , \R_DATA_TEMPR1[27] , 
        \R_DATA_TEMPR1[26] , \R_DATA_TEMPR1[25] , \R_DATA_TEMPR1[24] , 
        \R_DATA_TEMPR1[23] , \R_DATA_TEMPR1[22] , \R_DATA_TEMPR1[21] , 
        \R_DATA_TEMPR1[20] }));
    OR4 OR4_355 (.A(\R_DATA_TEMPR4[29] ), .B(\R_DATA_TEMPR5[29] ), .C(
        \R_DATA_TEMPR6[29] ), .D(\R_DATA_TEMPR7[29] ), .Y(OR4_355_Y));
    OR4 OR4_344 (.A(OR4_228_Y), .B(OR4_150_Y), .C(OR4_102_Y), .D(
        OR4_120_Y), .Y(OR4_344_Y));
    OR4 OR4_328 (.A(OR4_94_Y), .B(OR4_146_Y), .C(OR4_145_Y), .D(
        OR4_207_Y), .Y(OR4_328_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R13C0 (.BLK_EN(\BLKX0[13] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][0] ), .R_DATA({nc52, nc53, 
        \R_DATA_TEMPR13[9] , \R_DATA_TEMPR13[8] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR13[6] , \R_DATA_TEMPR13[5] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR13[3] , \R_DATA_TEMPR13[2] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR13[0] }));
    OR4 OR4_185 (.A(\R_DATA_TEMPR28[14] ), .B(\R_DATA_TEMPR29[14] ), 
        .C(\R_DATA_TEMPR30[14] ), .D(\R_DATA_TEMPR31[14] ), .Y(
        OR4_185_Y));
    OR4 OR4_141 (.A(\R_DATA_TEMPR24[20] ), .B(\R_DATA_TEMPR25[20] ), 
        .C(\R_DATA_TEMPR26[20] ), .D(\R_DATA_TEMPR27[20] ), .Y(
        OR4_141_Y));
    OR4 OR4_36 (.A(\R_DATA_TEMPR12[22] ), .B(\R_DATA_TEMPR13[22] ), .C(
        \R_DATA_TEMPR14[22] ), .D(\R_DATA_TEMPR15[22] ), .Y(OR4_36_Y));
    CFG3 #( .INIT(8'h40) )  CFG3_23 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_23_Y));
    OR4 OR4_21 (.A(\R_DATA_TEMPR16[23] ), .B(\R_DATA_TEMPR17[23] ), .C(
        \R_DATA_TEMPR18[23] ), .D(\R_DATA_TEMPR19[23] ), .Y(OR4_21_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[14]  (.A(CFG3_2_Y), .B(
        CFG3_17_Y), .Y(\BLKX0[14] ));
    OR4 OR4_129 (.A(OR4_349_Y), .B(OR2_7_Y), .C(\R_DATA_TEMPR22[15] ), 
        .D(\R_DATA_TEMPR23[15] ), .Y(OR4_129_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R20C1 (.BLK_EN(\BLKX0[20] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[20] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][1] ), .R_DATA({nc54, nc55, 
        \R_DATA_TEMPR20[19] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR20[17] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR20[15] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR20[13] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR20[11] , \R_DATA_TEMPR20[10] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[18]  (.A(CFG3_16_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[18] ));
    OR4 OR4_285 (.A(OR4_59_Y), .B(OR4_275_Y), .C(OR4_290_Y), .D(
        OR4_115_Y), .Y(OR4_285_Y));
    OR4 OR4_202 (.A(\R_DATA_TEMPR28[21] ), .B(\R_DATA_TEMPR29[21] ), 
        .C(\R_DATA_TEMPR30[21] ), .D(\R_DATA_TEMPR31[21] ), .Y(
        OR4_202_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_13 (.A(W_EN), .B(W_ADDR[10]), .C(
        W_ADDR[9]), .Y(CFG3_13_Y));
    OR4 OR4_272 (.A(\R_DATA_TEMPR4[30] ), .B(\R_DATA_TEMPR5[30] ), .C(
        \R_DATA_TEMPR6[30] ), .D(\R_DATA_TEMPR7[30] ), .Y(OR4_272_Y));
    OR4 OR4_44 (.A(\R_DATA_TEMPR4[7] ), .B(\R_DATA_TEMPR5[7] ), .C(
        \R_DATA_TEMPR6[7] ), .D(\R_DATA_TEMPR7[7] ), .Y(OR4_44_Y));
    OR4 OR4_300 (.A(\R_DATA_TEMPR12[14] ), .B(\R_DATA_TEMPR13[14] ), 
        .C(\R_DATA_TEMPR14[14] ), .D(\R_DATA_TEMPR15[14] ), .Y(
        OR4_300_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[31]  (.A(CFG3_15_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[31] ));
    OR4 OR4_288 (.A(\R_DATA_TEMPR4[5] ), .B(\R_DATA_TEMPR5[5] ), .C(
        \R_DATA_TEMPR6[5] ), .D(\R_DATA_TEMPR7[5] ), .Y(OR4_288_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_0 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_0_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R2C2 (.BLK_EN(\BLKX0[2] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][2] ), .R_DATA({nc56, nc57, 
        \R_DATA_TEMPR2[29] , \R_DATA_TEMPR2[28] , \R_DATA_TEMPR2[27] , 
        \R_DATA_TEMPR2[26] , \R_DATA_TEMPR2[25] , \R_DATA_TEMPR2[24] , 
        \R_DATA_TEMPR2[23] , \R_DATA_TEMPR2[22] , \R_DATA_TEMPR2[21] , 
        \R_DATA_TEMPR2[20] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[7]  (.A(CFG3_15_Y), .B(CFG3_5_Y)
        , .Y(\BLKX0[7] ));
    OR4 OR4_30 (.A(\R_DATA_TEMPR8[14] ), .B(\R_DATA_TEMPR9[14] ), .C(
        \R_DATA_TEMPR10[14] ), .D(\R_DATA_TEMPR11[14] ), .Y(OR4_30_Y));
    OR4 OR4_297 (.A(OR4_287_Y), .B(OR4_283_Y), .C(OR4_255_Y), .D(
        OR4_353_Y), .Y(OR4_297_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R13C3 (.BLK_EN(\BLKX0[13] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][3] ), .R_DATA({nc58, nc59, 
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR13[38] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR13[36] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR13[34] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR13[32] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR13[30] }));
    OR4 OR4_37 (.A(\R_DATA_TEMPR12[20] ), .B(\R_DATA_TEMPR13[20] ), .C(
        \R_DATA_TEMPR14[20] ), .D(\R_DATA_TEMPR15[20] ), .Y(OR4_37_Y));
    OR4 OR4_197 (.A(\R_DATA_TEMPR8[9] ), .B(\R_DATA_TEMPR9[9] ), .C(
        \R_DATA_TEMPR10[9] ), .D(\R_DATA_TEMPR11[9] ), .Y(OR4_197_Y));
    OR4 OR4_357 (.A(\R_DATA_TEMPR4[33] ), .B(\R_DATA_TEMPR5[33] ), .C(
        \R_DATA_TEMPR6[33] ), .D(\R_DATA_TEMPR7[33] ), .Y(OR4_357_Y));
    OR4 OR4_150 (.A(\R_DATA_TEMPR4[18] ), .B(\R_DATA_TEMPR5[18] ), .C(
        \R_DATA_TEMPR6[18] ), .D(\R_DATA_TEMPR7[18] ), .Y(OR4_150_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_20 (.A(W_EN), .B(W_ADDR[10]), .C(
        W_ADDR[9]), .Y(CFG3_20_Y));
    OR4 OR4_163 (.A(\R_DATA_TEMPR24[22] ), .B(\R_DATA_TEMPR25[22] ), 
        .C(\R_DATA_TEMPR26[22] ), .D(\R_DATA_TEMPR27[22] ), .Y(
        OR4_163_Y));
    OR4 OR4_343 (.A(OR4_50_Y), .B(OR2_5_Y), .C(\R_DATA_TEMPR22[5] ), 
        .D(\R_DATA_TEMPR23[5] ), .Y(OR4_343_Y));
    OR4 OR4_336 (.A(\R_DATA_TEMPR0[13] ), .B(\R_DATA_TEMPR1[13] ), .C(
        \R_DATA_TEMPR2[13] ), .D(\R_DATA_TEMPR3[13] ), .Y(OR4_336_Y));
    OR4 OR4_294 (.A(OR4_266_Y), .B(OR4_186_Y), .C(OR4_270_Y), .D(
        OR4_73_Y), .Y(OR4_294_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R29C1 (.BLK_EN(\BLKX0[29] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[29] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][1] ), .R_DATA({nc60, nc61, 
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR29[18] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR29[16] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR29[14] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR29[12] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR29[10] }));
    OR4 \OR4_R_DATA[24]  (.A(OR4_308_Y), .B(OR4_181_Y), .C(OR4_1_Y), 
        .D(OR4_152_Y), .Y(R_DATA[24]));
    OR4 OR4_85 (.A(\R_DATA_TEMPR12[28] ), .B(\R_DATA_TEMPR13[28] ), .C(
        \R_DATA_TEMPR14[28] ), .D(\R_DATA_TEMPR15[28] ), .Y(OR4_85_Y));
    OR4 OR4_146 (.A(\R_DATA_TEMPR4[21] ), .B(\R_DATA_TEMPR5[21] ), .C(
        \R_DATA_TEMPR6[21] ), .D(\R_DATA_TEMPR7[21] ), .Y(OR4_146_Y));
    OR4 OR4_158 (.A(\R_DATA_TEMPR4[6] ), .B(\R_DATA_TEMPR5[6] ), .C(
        \R_DATA_TEMPR6[6] ), .D(\R_DATA_TEMPR7[6] ), .Y(OR4_158_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_256_Y), .B(OR4_245_Y), .C(OR4_196_Y), 
        .D(OR4_29_Y), .Y(R_DATA[12]));
    CFG3 #( .INIT(8'h80) )  CFG3_10 (.A(W_EN), .B(W_ADDR[10]), .C(
        W_ADDR[9]), .Y(CFG3_10_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[29]  (.A(CFG3_12_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[29] ));
    OR4 OR4_69 (.A(\R_DATA_TEMPR16[6] ), .B(\R_DATA_TEMPR17[6] ), .C(
        \R_DATA_TEMPR18[6] ), .D(\R_DATA_TEMPR19[6] ), .Y(OR4_69_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[8]  (.A(CFG3_11_Y), .B(
        CFG3_20_Y), .Y(\BLKZ0[8] ));
    OR4 OR4_227 (.A(\R_DATA_TEMPR8[23] ), .B(\R_DATA_TEMPR9[23] ), .C(
        \R_DATA_TEMPR10[23] ), .D(\R_DATA_TEMPR11[23] ), .Y(OR4_227_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R5C2 (.BLK_EN(\BLKX0[5] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][2] ), .R_DATA({nc62, nc63, 
        \R_DATA_TEMPR5[29] , \R_DATA_TEMPR5[28] , \R_DATA_TEMPR5[27] , 
        \R_DATA_TEMPR5[26] , \R_DATA_TEMPR5[25] , \R_DATA_TEMPR5[24] , 
        \R_DATA_TEMPR5[23] , \R_DATA_TEMPR5[22] , \R_DATA_TEMPR5[21] , 
        \R_DATA_TEMPR5[20] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[25]  (.A(CFG3_1_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[25] ));
    OR4 OR4_127 (.A(\R_DATA_TEMPR0[11] ), .B(\R_DATA_TEMPR1[11] ), .C(
        \R_DATA_TEMPR2[11] ), .D(\R_DATA_TEMPR3[11] ), .Y(OR4_127_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[10]  (.A(CFG3_8_Y), .B(
        CFG3_17_Y), .Y(\BLKX0[10] ));
    OR4 OR4_348 (.A(\R_DATA_TEMPR8[33] ), .B(\R_DATA_TEMPR9[33] ), .C(
        \R_DATA_TEMPR10[33] ), .D(\R_DATA_TEMPR11[33] ), .Y(OR4_348_Y));
    OR4 OR4_162 (.A(\R_DATA_TEMPR28[36] ), .B(\R_DATA_TEMPR29[36] ), 
        .C(\R_DATA_TEMPR30[36] ), .D(\R_DATA_TEMPR31[36] ), .Y(
        OR4_162_Y));
    OR4 OR4_282 (.A(\R_DATA_TEMPR24[32] ), .B(\R_DATA_TEMPR25[32] ), 
        .C(\R_DATA_TEMPR26[32] ), .D(\R_DATA_TEMPR27[32] ), .Y(
        OR4_282_Y));
    OR4 OR4_316 (.A(\R_DATA_TEMPR8[3] ), .B(\R_DATA_TEMPR9[3] ), .C(
        \R_DATA_TEMPR10[3] ), .D(\R_DATA_TEMPR11[3] ), .Y(OR4_316_Y));
    OR4 OR4_134 (.A(\R_DATA_TEMPR24[8] ), .B(\R_DATA_TEMPR25[8] ), .C(
        \R_DATA_TEMPR26[8] ), .D(\R_DATA_TEMPR27[8] ), .Y(OR4_134_Y));
    OR2 OR2_35 (.A(\R_DATA_TEMPR20[0] ), .B(\R_DATA_TEMPR21[0] ), .Y(
        OR2_35_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R21C0 (.BLK_EN(\BLKX0[21] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[21] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][0] ), .R_DATA({nc64, nc65, 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR21[4] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR21[1] , 
        \R_DATA_TEMPR21[0] }));
    OR4 OR4_103 (.A(OR4_144_Y), .B(OR2_11_Y), .C(\R_DATA_TEMPR22[30] ), 
        .D(\R_DATA_TEMPR23[30] ), .Y(OR4_103_Y));
    OR4 OR4_224 (.A(\R_DATA_TEMPR24[7] ), .B(\R_DATA_TEMPR25[7] ), .C(
        \R_DATA_TEMPR26[7] ), .D(\R_DATA_TEMPR27[7] ), .Y(OR4_224_Y));
    OR4 OR4_149 (.A(\R_DATA_TEMPR28[4] ), .B(\R_DATA_TEMPR29[4] ), .C(
        \R_DATA_TEMPR30[4] ), .D(\R_DATA_TEMPR31[4] ), .Y(OR4_149_Y));
    OR4 \OR4_R_DATA[13]  (.A(OR4_212_Y), .B(OR4_130_Y), .C(OR4_114_Y), 
        .D(OR4_106_Y), .Y(R_DATA[13]));
    OR4 OR4_173 (.A(\R_DATA_TEMPR28[18] ), .B(\R_DATA_TEMPR29[18] ), 
        .C(\R_DATA_TEMPR30[18] ), .D(\R_DATA_TEMPR31[18] ), .Y(
        OR4_173_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R0C0 (.BLK_EN(\BLKX0[0] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][0] ), .R_DATA({nc66, nc67, 
        \R_DATA_TEMPR0[9] , \R_DATA_TEMPR0[8] , \R_DATA_TEMPR0[7] , 
        \R_DATA_TEMPR0[6] , \R_DATA_TEMPR0[5] , \R_DATA_TEMPR0[4] , 
        \R_DATA_TEMPR0[3] , \R_DATA_TEMPR0[2] , \R_DATA_TEMPR0[1] , 
        \R_DATA_TEMPR0[0] }));
    OR4 OR4_269 (.A(\R_DATA_TEMPR28[8] ), .B(\R_DATA_TEMPR29[8] ), .C(
        \R_DATA_TEMPR30[8] ), .D(\R_DATA_TEMPR31[8] ), .Y(OR4_269_Y));
    OR4 OR4_62 (.A(\R_DATA_TEMPR16[22] ), .B(\R_DATA_TEMPR17[22] ), .C(
        \R_DATA_TEMPR18[22] ), .D(\R_DATA_TEMPR19[22] ), .Y(OR4_62_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R2C1 (.BLK_EN(\BLKX0[2] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][1] ), .R_DATA({nc68, nc69, 
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR2[18] , \R_DATA_TEMPR2[17] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR2[15] , \R_DATA_TEMPR2[14] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR2[12] , \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR2[10] }));
    OR4 OR4_38 (.A(\R_DATA_TEMPR12[39] ), .B(\R_DATA_TEMPR13[39] ), .C(
        \R_DATA_TEMPR14[39] ), .D(\R_DATA_TEMPR15[39] ), .Y(OR4_38_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R3C0 (.BLK_EN(\BLKX0[3] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][0] ), .R_DATA({nc70, nc71, 
        \R_DATA_TEMPR3[9] , \R_DATA_TEMPR3[8] , \R_DATA_TEMPR3[7] , 
        \R_DATA_TEMPR3[6] , \R_DATA_TEMPR3[5] , \R_DATA_TEMPR3[4] , 
        \R_DATA_TEMPR3[3] , \R_DATA_TEMPR3[2] , \R_DATA_TEMPR3[1] , 
        \R_DATA_TEMPR3[0] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[18]  (.A(CFG3_8_Y), .B(CFG3_9_Y)
        , .Y(\BLKX0[18] ));
    OR4 OR4_325 (.A(OR4_101_Y), .B(OR2_25_Y), .C(\R_DATA_TEMPR22[7] ), 
        .D(\R_DATA_TEMPR23[7] ), .Y(OR4_325_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R20C3 (.BLK_EN(\BLKX0[20] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[20] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][3] ), .R_DATA({nc72, nc73, 
        \R_DATA_TEMPR20[39] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR20[37] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR20[35] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR20[33] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR20[31] , \R_DATA_TEMPR20[30] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[13]  (.A(CFG3_12_Y), .B(
        CFG3_17_Y), .Y(\BLKX0[13] ));
    OR4 OR4_114 (.A(\R_DATA_TEMPR24[13] ), .B(\R_DATA_TEMPR25[13] ), 
        .C(\R_DATA_TEMPR26[13] ), .D(\R_DATA_TEMPR27[13] ), .Y(
        OR4_114_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[0]  (.A(CFG3_11_Y), .B(CFG3_4_Y)
        , .Y(\BLKZ0[0] ));
    OR4 OR4_155 (.A(\R_DATA_TEMPR16[29] ), .B(\R_DATA_TEMPR17[29] ), 
        .C(\R_DATA_TEMPR18[29] ), .D(\R_DATA_TEMPR19[29] ), .Y(
        OR4_155_Y));
    OR4 OR4_102 (.A(\R_DATA_TEMPR8[18] ), .B(\R_DATA_TEMPR9[18] ), .C(
        \R_DATA_TEMPR10[18] ), .D(\R_DATA_TEMPR11[18] ), .Y(OR4_102_Y));
    OR4 OR4_172 (.A(\R_DATA_TEMPR16[32] ), .B(\R_DATA_TEMPR17[32] ), 
        .C(\R_DATA_TEMPR18[32] ), .D(\R_DATA_TEMPR19[32] ), .Y(
        OR4_172_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R16C0 (.BLK_EN(\BLKX0[16] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][0] ), .R_DATA({nc74, nc75, 
        \R_DATA_TEMPR16[9] , \R_DATA_TEMPR16[8] , \R_DATA_TEMPR16[7] , 
        \R_DATA_TEMPR16[6] , \R_DATA_TEMPR16[5] , \R_DATA_TEMPR16[4] , 
        \R_DATA_TEMPR16[3] , \R_DATA_TEMPR16[2] , \R_DATA_TEMPR16[1] , 
        \R_DATA_TEMPR16[0] }));
    OR4 OR4_255 (.A(\R_DATA_TEMPR8[0] ), .B(\R_DATA_TEMPR9[0] ), .C(
        \R_DATA_TEMPR10[0] ), .D(\R_DATA_TEMPR11[0] ), .Y(OR4_255_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R8C0 (.BLK_EN(\BLKX0[8] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][0] ), .R_DATA({nc76, nc77, 
        \R_DATA_TEMPR8[9] , \R_DATA_TEMPR8[8] , \R_DATA_TEMPR8[7] , 
        \R_DATA_TEMPR8[6] , \R_DATA_TEMPR8[5] , \R_DATA_TEMPR8[4] , 
        \R_DATA_TEMPR8[3] , \R_DATA_TEMPR8[2] , \R_DATA_TEMPR8[1] , 
        \R_DATA_TEMPR8[0] }));
    OR4 OR4_190 (.A(\R_DATA_TEMPR8[8] ), .B(\R_DATA_TEMPR9[8] ), .C(
        \R_DATA_TEMPR10[8] ), .D(\R_DATA_TEMPR11[8] ), .Y(OR4_190_Y));
    OR4 OR4_26 (.A(OR4_189_Y), .B(OR2_28_Y), .C(\R_DATA_TEMPR22[19] ), 
        .D(\R_DATA_TEMPR23[19] ), .Y(OR4_26_Y));
    OR4 OR4_53 (.A(\R_DATA_TEMPR16[13] ), .B(\R_DATA_TEMPR17[13] ), .C(
        \R_DATA_TEMPR18[13] ), .D(\R_DATA_TEMPR19[13] ), .Y(OR4_53_Y));
    OR4 OR4_209 (.A(\R_DATA_TEMPR16[1] ), .B(\R_DATA_TEMPR17[1] ), .C(
        \R_DATA_TEMPR18[1] ), .D(\R_DATA_TEMPR19[1] ), .Y(OR4_209_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R3C3 (.BLK_EN(\BLKX0[3] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][3] ), .R_DATA({nc78, nc79, 
        \R_DATA_TEMPR3[39] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR3[37] , 
        \R_DATA_TEMPR3[36] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR3[34] , 
        \R_DATA_TEMPR3[33] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR3[31] , 
        \R_DATA_TEMPR3[30] }));
    OR4 OR4_279 (.A(\R_DATA_TEMPR28[9] ), .B(\R_DATA_TEMPR29[9] ), .C(
        \R_DATA_TEMPR30[9] ), .D(\R_DATA_TEMPR31[9] ), .Y(OR4_279_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R30C1 (.BLK_EN(\BLKX0[30] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[30] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][1] ), .R_DATA({nc80, nc81, 
        \R_DATA_TEMPR30[19] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR30[17] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR30[15] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR30[13] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR30[11] , \R_DATA_TEMPR30[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R18C0 (.BLK_EN(\BLKX0[18] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][0] ), .R_DATA({nc82, nc83, 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR18[7] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR18[4] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR18[1] , 
        \R_DATA_TEMPR18[0] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[12]  (.A(CFG3_18_Y), .B(
        CFG3_20_Y), .Y(\BLKZ0[12] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[24]  (.A(CFG3_11_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[24] ));
    OR4 OR4_89 (.A(OR4_110_Y), .B(OR4_221_Y), .C(OR4_316_Y), .D(
        OR4_123_Y), .Y(OR4_89_Y));
    OR4 OR4_198 (.A(\R_DATA_TEMPR0[28] ), .B(\R_DATA_TEMPR1[28] ), .C(
        \R_DATA_TEMPR2[28] ), .D(\R_DATA_TEMPR3[28] ), .Y(OR4_198_Y));
    OR4 OR4_258 (.A(\R_DATA_TEMPR8[13] ), .B(\R_DATA_TEMPR9[13] ), .C(
        \R_DATA_TEMPR10[13] ), .D(\R_DATA_TEMPR11[13] ), .Y(OR4_258_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_328_Y), .B(OR4_311_Y), .C(OR4_320_Y), 
        .D(OR4_202_Y), .Y(R_DATA[21]));
    OR4 OR4_183 (.A(\R_DATA_TEMPR16[38] ), .B(\R_DATA_TEMPR17[38] ), 
        .C(\R_DATA_TEMPR18[38] ), .D(\R_DATA_TEMPR19[38] ), .Y(
        OR4_183_Y));
    OR4 OR4_332 (.A(\R_DATA_TEMPR8[32] ), .B(\R_DATA_TEMPR9[32] ), .C(
        \R_DATA_TEMPR10[32] ), .D(\R_DATA_TEMPR11[32] ), .Y(OR4_332_Y));
    OR4 OR4_13 (.A(OR4_67_Y), .B(OR2_4_Y), .C(\R_DATA_TEMPR22[10] ), 
        .D(\R_DATA_TEMPR23[10] ), .Y(OR4_13_Y));
    OR4 OR4_247 (.A(\R_DATA_TEMPR8[12] ), .B(\R_DATA_TEMPR9[12] ), .C(
        \R_DATA_TEMPR10[12] ), .D(\R_DATA_TEMPR11[12] ), .Y(OR4_247_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R9C2 (.BLK_EN(\BLKX0[9] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][2] ), .R_DATA({nc84, nc85, 
        \R_DATA_TEMPR9[29] , \R_DATA_TEMPR9[28] , \R_DATA_TEMPR9[27] , 
        \R_DATA_TEMPR9[26] , \R_DATA_TEMPR9[25] , \R_DATA_TEMPR9[24] , 
        \R_DATA_TEMPR9[23] , \R_DATA_TEMPR9[22] , \R_DATA_TEMPR9[21] , 
        \R_DATA_TEMPR9[20] }));
    CFG3 #( .INIT(8'h80) )  CFG3_3 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_3_Y));
    OR4 OR4_327 (.A(\R_DATA_TEMPR4[24] ), .B(\R_DATA_TEMPR5[24] ), .C(
        \R_DATA_TEMPR6[24] ), .D(\R_DATA_TEMPR7[24] ), .Y(OR4_327_Y));
    OR4 OR4_147 (.A(\R_DATA_TEMPR12[32] ), .B(\R_DATA_TEMPR13[32] ), 
        .C(\R_DATA_TEMPR14[32] ), .D(\R_DATA_TEMPR15[32] ), .Y(
        OR4_147_Y));
    OR4 OR4_120 (.A(\R_DATA_TEMPR12[18] ), .B(\R_DATA_TEMPR13[18] ), 
        .C(\R_DATA_TEMPR14[18] ), .D(\R_DATA_TEMPR15[18] ), .Y(
        OR4_120_Y));
    OR4 OR4_51 (.A(OR4_157_Y), .B(OR4_288_Y), .C(OR4_252_Y), .D(
        OR4_112_Y), .Y(OR4_51_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[6]  (.A(CFG3_7_Y), .B(CFG3_4_Y), 
        .Y(\BLKZ0[6] ));
    OR2 OR2_2 (.A(\R_DATA_TEMPR20[26] ), .B(\R_DATA_TEMPR21[26] ), .Y(
        OR2_2_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[21]  (.A(CFG3_12_Y), .B(
        CFG3_9_Y), .Y(\BLKX0[21] ));
    OR4 \OR4_R_DATA[20]  (.A(OR4_262_Y), .B(OR4_351_Y), .C(OR4_141_Y), 
        .D(OR4_10_Y), .Y(R_DATA[20]));
    OR2 OR2_39 (.A(\R_DATA_TEMPR20[29] ), .B(\R_DATA_TEMPR21[29] ), .Y(
        OR2_39_Y));
    OR4 OR4_20 (.A(\R_DATA_TEMPR16[4] ), .B(\R_DATA_TEMPR17[4] ), .C(
        \R_DATA_TEMPR18[4] ), .D(\R_DATA_TEMPR19[4] ), .Y(OR4_20_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[19]  (.A(CFG3_23_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[19] ));
    OR4 \OR4_R_DATA[26]  (.A(OR4_135_Y), .B(OR4_331_Y), .C(OR4_28_Y), 
        .D(OR4_48_Y), .Y(R_DATA[26]));
    OR4 OR4_244 (.A(OR4_195_Y), .B(OR2_24_Y), .C(\R_DATA_TEMPR22[17] ), 
        .D(\R_DATA_TEMPR23[17] ), .Y(OR4_244_Y));
    OR4 OR4_27 (.A(OR4_168_Y), .B(OR4_18_Y), .C(OR4_34_Y), .D(
        OR4_218_Y), .Y(OR4_27_Y));
    OR4 OR4_82 (.A(OR4_43_Y), .B(OR4_158_Y), .C(OR4_90_Y), .D(OR4_87_Y)
        , .Y(OR4_82_Y));
    OR4 OR4_128 (.A(\R_DATA_TEMPR28[30] ), .B(\R_DATA_TEMPR29[30] ), 
        .C(\R_DATA_TEMPR30[30] ), .D(\R_DATA_TEMPR31[30] ), .Y(
        OR4_128_Y));
    OR4 OR4_230 (.A(\R_DATA_TEMPR24[25] ), .B(\R_DATA_TEMPR25[25] ), 
        .C(\R_DATA_TEMPR26[25] ), .D(\R_DATA_TEMPR27[25] ), .Y(
        OR4_230_Y));
    OR4 OR4_182 (.A(\R_DATA_TEMPR16[9] ), .B(\R_DATA_TEMPR17[9] ), .C(
        \R_DATA_TEMPR18[9] ), .D(\R_DATA_TEMPR19[9] ), .Y(OR4_182_Y));
    OR4 OR4_312 (.A(OR4_96_Y), .B(OR4_302_Y), .C(OR4_319_Y), .D(
        OR4_136_Y), .Y(OR4_312_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R24C3 (.BLK_EN(\BLKX0[24] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[24] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][3] ), .R_DATA({nc86, nc87, 
        \R_DATA_TEMPR24[39] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR24[37] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR24[35] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR24[33] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR24[31] , \R_DATA_TEMPR24[30] }));
    OR4 OR4_64 (.A(\R_DATA_TEMPR16[35] ), .B(\R_DATA_TEMPR17[35] ), .C(
        \R_DATA_TEMPR18[35] ), .D(\R_DATA_TEMPR19[35] ), .Y(OR4_64_Y));
    OR4 OR4_11 (.A(\R_DATA_TEMPR24[6] ), .B(\R_DATA_TEMPR25[6] ), .C(
        \R_DATA_TEMPR26[6] ), .D(\R_DATA_TEMPR27[6] ), .Y(OR4_11_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R24C1 (.BLK_EN(\BLKX0[24] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[24] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][1] ), .R_DATA({nc88, nc89, 
        \R_DATA_TEMPR24[19] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR24[17] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR24[15] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR24[13] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR24[11] , \R_DATA_TEMPR24[10] }));
    OR4 OR4_345 (.A(OR4_42_Y), .B(OR4_257_Y), .C(OR4_332_Y), .D(
        OR4_147_Y), .Y(OR4_345_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R1C3 (.BLK_EN(\BLKX0[1] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][3] ), .R_DATA({nc90, nc91, 
        \R_DATA_TEMPR1[39] , \R_DATA_TEMPR1[38] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR1[36] , \R_DATA_TEMPR1[35] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR1[33] , \R_DATA_TEMPR1[32] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR1[30] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R27C2 (.BLK_EN(\BLKX0[27] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[27] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][2] ), .R_DATA({nc92, nc93, 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR27[28] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR27[26] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR27[24] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR27[22] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR27[20] }));
    OR4 OR4_236 (.A(\R_DATA_TEMPR24[1] ), .B(\R_DATA_TEMPR25[1] ), .C(
        \R_DATA_TEMPR26[1] ), .D(\R_DATA_TEMPR27[1] ), .Y(OR4_236_Y));
    OR2 OR2_7 (.A(\R_DATA_TEMPR20[15] ), .B(\R_DATA_TEMPR21[15] ), .Y(
        OR2_7_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R17C3 (.BLK_EN(\BLKX0[17] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][3] ), .R_DATA({nc94, nc95, 
        \R_DATA_TEMPR17[39] , \R_DATA_TEMPR17[38] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR17[36] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR17[34] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR17[32] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR17[30] }));
    OR4 OR4_73 (.A(\R_DATA_TEMPR12[10] ), .B(\R_DATA_TEMPR13[10] ), .C(
        \R_DATA_TEMPR14[10] ), .D(\R_DATA_TEMPR15[10] ), .Y(OR4_73_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[17]  (.A(CFG3_1_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[17] ));
    OR4 OR4_195 (.A(\R_DATA_TEMPR16[17] ), .B(\R_DATA_TEMPR17[17] ), 
        .C(\R_DATA_TEMPR18[17] ), .D(\R_DATA_TEMPR19[17] ), .Y(
        OR4_195_Y));
    OR4 OR4_252 (.A(\R_DATA_TEMPR8[5] ), .B(\R_DATA_TEMPR9[5] ), .C(
        \R_DATA_TEMPR10[5] ), .D(\R_DATA_TEMPR11[5] ), .Y(OR4_252_Y));
    OR4 OR4_289 (.A(\R_DATA_TEMPR12[26] ), .B(\R_DATA_TEMPR13[26] ), 
        .C(\R_DATA_TEMPR14[26] ), .D(\R_DATA_TEMPR15[26] ), .Y(
        OR4_289_Y));
    OR2 OR2_32 (.A(\R_DATA_TEMPR20[39] ), .B(\R_DATA_TEMPR21[39] ), .Y(
        OR2_32_Y));
    OR2 OR2_1 (.A(\R_DATA_TEMPR20[33] ), .B(\R_DATA_TEMPR21[33] ), .Y(
        OR2_1_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R19C0 (.BLK_EN(\BLKX0[19] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][0] ), .R_DATA({nc96, nc97, 
        \R_DATA_TEMPR19[9] , \R_DATA_TEMPR19[8] , \R_DATA_TEMPR19[7] , 
        \R_DATA_TEMPR19[6] , \R_DATA_TEMPR19[5] , \R_DATA_TEMPR19[4] , 
        \R_DATA_TEMPR19[3] , \R_DATA_TEMPR19[2] , \R_DATA_TEMPR19[1] , 
        \R_DATA_TEMPR19[0] }));
    OR4 OR4_210 (.A(OR4_309_Y), .B(OR2_12_Y), .C(\R_DATA_TEMPR22[14] ), 
        .D(\R_DATA_TEMPR23[14] ), .Y(OR4_210_Y));
    OR4 OR4_350 (.A(\R_DATA_TEMPR0[7] ), .B(\R_DATA_TEMPR1[7] ), .C(
        \R_DATA_TEMPR2[7] ), .D(\R_DATA_TEMPR3[7] ), .Y(OR4_350_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R0C3 (.BLK_EN(\BLKX0[0] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][3] ), .R_DATA({nc98, nc99, 
        \R_DATA_TEMPR0[39] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR0[37] , 
        \R_DATA_TEMPR0[36] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR0[34] , 
        \R_DATA_TEMPR0[33] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR0[31] , 
        \R_DATA_TEMPR0[30] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[5]  (.A(CFG3_12_Y), .B(CFG3_5_Y)
        , .Y(\BLKX0[5] ));
    OR4 OR4_295 (.A(OR4_108_Y), .B(OR2_13_Y), .C(\R_DATA_TEMPR22[18] ), 
        .D(\R_DATA_TEMPR23[18] ), .Y(OR4_295_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R19C3 (.BLK_EN(\BLKX0[19] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][3] ), .R_DATA({nc100, nc101, 
        \R_DATA_TEMPR19[39] , \R_DATA_TEMPR19[38] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR19[36] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR19[34] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR19[32] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR19[30] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R25C1 (.BLK_EN(\BLKX0[25] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[25] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][1] ), .R_DATA({nc102, nc103, 
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR25[18] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR25[16] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR25[14] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR25[12] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR25[10] }));
    OR4 OR4_35 (.A(\R_DATA_TEMPR0[4] ), .B(\R_DATA_TEMPR1[4] ), .C(
        \R_DATA_TEMPR2[4] ), .D(\R_DATA_TEMPR3[4] ), .Y(OR4_35_Y));
    OR4 OR4_216 (.A(\R_DATA_TEMPR8[22] ), .B(\R_DATA_TEMPR9[22] ), .C(
        \R_DATA_TEMPR10[22] ), .D(\R_DATA_TEMPR11[22] ), .Y(OR4_216_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R31C0 (.BLK_EN(\BLKX0[31] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[31] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][0] ), .R_DATA({nc104, nc105, 
        \R_DATA_TEMPR31[9] , \R_DATA_TEMPR31[8] , \R_DATA_TEMPR31[7] , 
        \R_DATA_TEMPR31[6] , \R_DATA_TEMPR31[5] , \R_DATA_TEMPR31[4] , 
        \R_DATA_TEMPR31[3] , \R_DATA_TEMPR31[2] , \R_DATA_TEMPR31[1] , 
        \R_DATA_TEMPR31[0] }));
    OR4 OR4_71 (.A(\R_DATA_TEMPR12[8] ), .B(\R_DATA_TEMPR13[8] ), .C(
        \R_DATA_TEMPR14[8] ), .D(\R_DATA_TEMPR15[8] ), .Y(OR4_71_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[9]  (.A(CFG3_1_Y), .B(CFG3_20_Y)
        , .Y(\BLKZ0[9] ));
    OR4 OR4_125 (.A(\R_DATA_TEMPR8[34] ), .B(\R_DATA_TEMPR9[34] ), .C(
        \R_DATA_TEMPR10[34] ), .D(\R_DATA_TEMPR11[34] ), .Y(OR4_125_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R20C0 (.BLK_EN(\BLKX0[20] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[20] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][0] ), .R_DATA({nc106, nc107, 
        \R_DATA_TEMPR20[9] , \R_DATA_TEMPR20[8] , \R_DATA_TEMPR20[7] , 
        \R_DATA_TEMPR20[6] , \R_DATA_TEMPR20[5] , \R_DATA_TEMPR20[4] , 
        \R_DATA_TEMPR20[3] , \R_DATA_TEMPR20[2] , \R_DATA_TEMPR20[1] , 
        \R_DATA_TEMPR20[0] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R21C3 (.BLK_EN(\BLKX0[21] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[21] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][3] ), .R_DATA({nc108, nc109, 
        \R_DATA_TEMPR21[39] , \R_DATA_TEMPR21[38] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR21[36] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR21[34] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR21[32] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR21[30] }));
    OR4 OR4_298 (.A(\R_DATA_TEMPR28[5] ), .B(\R_DATA_TEMPR29[5] ), .C(
        \R_DATA_TEMPR30[5] ), .D(\R_DATA_TEMPR31[5] ), .Y(OR4_298_Y));
    OR4 \OR4_R_DATA[27]  (.A(OR4_40_Y), .B(OR4_211_Y), .C(OR4_306_Y), 
        .D(OR4_347_Y), .Y(R_DATA[27]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R1C1 (.BLK_EN(\BLKX0[1] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][1] ), .R_DATA({nc110, nc111, 
        \R_DATA_TEMPR1[19] , \R_DATA_TEMPR1[18] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR1[16] , \R_DATA_TEMPR1[15] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR1[13] , \R_DATA_TEMPR1[12] , \R_DATA_TEMPR1[11] , 
        \R_DATA_TEMPR1[10] }));
    OR4 OR4_28 (.A(\R_DATA_TEMPR24[26] ), .B(\R_DATA_TEMPR25[26] ), .C(
        \R_DATA_TEMPR26[26] ), .D(\R_DATA_TEMPR27[26] ), .Y(OR4_28_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R30C3 (.BLK_EN(\BLKX0[30] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[30] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][3] ), .R_DATA({nc112, nc113, 
        \R_DATA_TEMPR30[39] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR30[37] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR30[35] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR30[33] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR30[31] , \R_DATA_TEMPR30[30] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R10C1 (.BLK_EN(\BLKX0[10] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][1] ), .R_DATA({nc114, nc115, 
        \R_DATA_TEMPR10[19] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR10[17] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR10[15] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR10[13] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR10[11] , \R_DATA_TEMPR10[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R26C3 (.BLK_EN(\BLKX0[26] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[26] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][3] ), .R_DATA({nc116, nc117, 
        \R_DATA_TEMPR26[39] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR26[37] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR26[35] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR26[33] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR26[31] , \R_DATA_TEMPR26[30] }));
    OR4 OR4_164 (.A(\R_DATA_TEMPR16[36] ), .B(\R_DATA_TEMPR17[36] ), 
        .C(\R_DATA_TEMPR18[36] ), .D(\R_DATA_TEMPR19[36] ), .Y(
        OR4_164_Y));
    OR4 OR4_225 (.A(OR4_296_Y), .B(OR4_140_Y), .C(OR4_216_Y), .D(
        OR4_36_Y), .Y(OR4_225_Y));
    OR4 OR4_347 (.A(\R_DATA_TEMPR28[27] ), .B(\R_DATA_TEMPR29[27] ), 
        .C(\R_DATA_TEMPR30[27] ), .D(\R_DATA_TEMPR31[27] ), .Y(
        OR4_347_Y));
    OR4 OR4_140 (.A(\R_DATA_TEMPR4[22] ), .B(\R_DATA_TEMPR5[22] ), .C(
        \R_DATA_TEMPR6[22] ), .D(\R_DATA_TEMPR7[22] ), .Y(OR4_140_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R23C2 (.BLK_EN(\BLKX0[23] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[23] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][2] ), .R_DATA({nc118, nc119, 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR23[28] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR23[26] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR23[24] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR23[22] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR23[20] }));
    OR4 OR4_306 (.A(\R_DATA_TEMPR24[27] ), .B(\R_DATA_TEMPR25[27] ), 
        .C(\R_DATA_TEMPR26[27] ), .D(\R_DATA_TEMPR27[27] ), .Y(
        OR4_306_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R6C1 (.BLK_EN(\BLKX0[6] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][1] ), .R_DATA({nc120, nc121, 
        \R_DATA_TEMPR6[19] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR6[17] , 
        \R_DATA_TEMPR6[16] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR6[14] , 
        \R_DATA_TEMPR6[13] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR6[11] , 
        \R_DATA_TEMPR6[10] }));
    OR4 OR4_84 (.A(OR4_223_Y), .B(OR4_355_Y), .C(OR4_138_Y), .D(
        OR4_291_Y), .Y(OR4_84_Y));
    OR4 OR4_148 (.A(\R_DATA_TEMPR12[30] ), .B(\R_DATA_TEMPR13[30] ), 
        .C(\R_DATA_TEMPR14[30] ), .D(\R_DATA_TEMPR15[30] ), .Y(
        OR4_148_Y));
    OR4 OR4_228 (.A(\R_DATA_TEMPR0[18] ), .B(\R_DATA_TEMPR1[18] ), .C(
        \R_DATA_TEMPR2[18] ), .D(\R_DATA_TEMPR3[18] ), .Y(OR4_228_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_4 (.A(W_EN), .B(W_ADDR[10]), .C(
        W_ADDR[9]), .Y(CFG3_4_Y));
    OR4 OR4_153 (.A(OR4_184_Y), .B(OR4_19_Y), .C(OR4_159_Y), .D(
        OR4_335_Y), .Y(OR4_153_Y));
    OR4 OR4_9 (.A(\R_DATA_TEMPR24[19] ), .B(\R_DATA_TEMPR25[19] ), .C(
        \R_DATA_TEMPR26[19] ), .D(\R_DATA_TEMPR27[19] ), .Y(OR4_9_Y));
    OR4 OR4_231 (.A(\R_DATA_TEMPR0[2] ), .B(\R_DATA_TEMPR1[2] ), .C(
        \R_DATA_TEMPR2[2] ), .D(\R_DATA_TEMPR3[2] ), .Y(OR4_231_Y));
    OR4 OR4_104 (.A(\R_DATA_TEMPR12[2] ), .B(\R_DATA_TEMPR13[2] ), .C(
        \R_DATA_TEMPR14[2] ), .D(\R_DATA_TEMPR15[2] ), .Y(OR4_104_Y));
    OR4 OR4_292 (.A(OR4_326_Y), .B(OR4_4_Y), .C(OR4_24_Y), .D(OR4_6_Y), 
        .Y(OR4_292_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_5 (.A(BLK_EN), .B(R_ADDR[10]), .C(
        R_ADDR[9]), .Y(CFG3_5_Y));
    OR4 OR4_174 (.A(OR4_47_Y), .B(OR4_75_Y), .C(OR4_190_Y), .D(
        OR4_71_Y), .Y(OR4_174_Y));
    OR2 OR2_34 (.A(\R_DATA_TEMPR20[1] ), .B(\R_DATA_TEMPR21[1] ), .Y(
        OR2_34_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[16]  (.A(CFG3_6_Y), .B(CFG3_9_Y)
        , .Y(\BLKX0[16] ));
    OR4 OR4_56 (.A(\R_DATA_TEMPR24[37] ), .B(\R_DATA_TEMPR25[37] ), .C(
        \R_DATA_TEMPR26[37] ), .D(\R_DATA_TEMPR27[37] ), .Y(OR4_56_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R19C1 (.BLK_EN(\BLKX0[19] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][1] ), .R_DATA({nc122, nc123, 
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR19[18] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR19[16] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR19[14] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR19[12] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR19[10] }));
    OR4 \OR4_R_DATA[2]  (.A(OR4_192_Y), .B(OR4_170_Y), .C(OR4_243_Y), 
        .D(OR4_274_Y), .Y(R_DATA[2]));
    OR4 OR4_152 (.A(\R_DATA_TEMPR28[24] ), .B(\R_DATA_TEMPR29[24] ), 
        .C(\R_DATA_TEMPR30[24] ), .D(\R_DATA_TEMPR31[24] ), .Y(
        OR4_152_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R25C3 (.BLK_EN(\BLKX0[25] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[25] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][3] ), .R_DATA({nc124, nc125, 
        \R_DATA_TEMPR25[39] , \R_DATA_TEMPR25[38] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR25[36] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR25[34] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR25[32] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR25[30] }));
    OR4 OR4_39 (.A(\R_DATA_TEMPR8[4] ), .B(\R_DATA_TEMPR9[4] ), .C(
        \R_DATA_TEMPR10[4] ), .D(\R_DATA_TEMPR11[4] ), .Y(OR4_39_Y));
    OR4 OR4_211 (.A(OR4_161_Y), .B(OR2_36_Y), .C(\R_DATA_TEMPR22[27] ), 
        .D(\R_DATA_TEMPR23[27] ), .Y(OR4_211_Y));
    OR2 OR2_9 (.A(\R_DATA_TEMPR20[3] ), .B(\R_DATA_TEMPR21[3] ), .Y(
        OR2_9_Y));
    OR4 OR4_145 (.A(\R_DATA_TEMPR8[21] ), .B(\R_DATA_TEMPR9[21] ), .C(
        \R_DATA_TEMPR10[21] ), .D(\R_DATA_TEMPR11[21] ), .Y(OR4_145_Y));
    OR4 OR4_222 (.A(\R_DATA_TEMPR24[5] ), .B(\R_DATA_TEMPR25[5] ), .C(
        \R_DATA_TEMPR26[5] ), .D(\R_DATA_TEMPR27[5] ), .Y(OR4_222_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R3C1 (.BLK_EN(\BLKX0[3] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[3] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][1] ), .R_DATA({nc126, nc127, 
        \R_DATA_TEMPR3[19] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR3[17] , 
        \R_DATA_TEMPR3[16] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR3[14] , 
        \R_DATA_TEMPR3[13] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR3[11] , 
        \R_DATA_TEMPR3[10] }));
    OR4 OR4_16 (.A(\R_DATA_TEMPR4[19] ), .B(\R_DATA_TEMPR5[19] ), .C(
        \R_DATA_TEMPR6[19] ), .D(\R_DATA_TEMPR7[19] ), .Y(OR4_16_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R9C0 (.BLK_EN(\BLKX0[9] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][0] ), .R_DATA({nc128, nc129, 
        \R_DATA_TEMPR9[9] , \R_DATA_TEMPR9[8] , \R_DATA_TEMPR9[7] , 
        \R_DATA_TEMPR9[6] , \R_DATA_TEMPR9[5] , \R_DATA_TEMPR9[4] , 
        \R_DATA_TEMPR9[3] , \R_DATA_TEMPR9[2] , \R_DATA_TEMPR9[1] , 
        \R_DATA_TEMPR9[0] }));
    OR4 OR4_259 (.A(\R_DATA_TEMPR24[30] ), .B(\R_DATA_TEMPR25[30] ), 
        .C(\R_DATA_TEMPR26[30] ), .D(\R_DATA_TEMPR27[30] ), .Y(
        OR4_259_Y));
    OR4 OR4_331 (.A(OR4_49_Y), .B(OR2_2_Y), .C(\R_DATA_TEMPR22[26] ), 
        .D(\R_DATA_TEMPR23[26] ), .Y(OR4_331_Y));
    OR4 OR4_4 (.A(\R_DATA_TEMPR4[1] ), .B(\R_DATA_TEMPR5[1] ), .C(
        \R_DATA_TEMPR6[1] ), .D(\R_DATA_TEMPR7[1] ), .Y(OR4_4_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[30]  (.A(CFG3_7_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[30] ));
    OR4 OR4_320 (.A(\R_DATA_TEMPR24[21] ), .B(\R_DATA_TEMPR25[21] ), 
        .C(\R_DATA_TEMPR26[21] ), .D(\R_DATA_TEMPR27[21] ), .Y(
        OR4_320_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R23C1 (.BLK_EN(\BLKX0[23] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[23] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][1] ), .R_DATA({nc130, nc131, 
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR23[18] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR23[16] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR23[14] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR23[12] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR23[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R11C0 (.BLK_EN(\BLKX0[11] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][0] ), .R_DATA({nc132, nc133, 
        \R_DATA_TEMPR11[9] , \R_DATA_TEMPR11[8] , \R_DATA_TEMPR11[7] , 
        \R_DATA_TEMPR11[6] , \R_DATA_TEMPR11[5] , \R_DATA_TEMPR11[4] , 
        \R_DATA_TEMPR11[3] , \R_DATA_TEMPR11[2] , \R_DATA_TEMPR11[1] , 
        \R_DATA_TEMPR11[0] }));
    OR4 \OR4_R_DATA[14]  (.A(OR4_342_Y), .B(OR4_210_Y), .C(OR4_23_Y), 
        .D(OR4_185_Y), .Y(R_DATA[14]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R27C0 (.BLK_EN(\BLKX0[27] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[27] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][0] ), .R_DATA({nc134, nc135, 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR27[7] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR27[4] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR27[0] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R22C0 (.BLK_EN(\BLKX0[22] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[22] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][0] ), .R_DATA({nc136, nc137, 
        \R_DATA_TEMPR22[9] , \R_DATA_TEMPR22[8] , \R_DATA_TEMPR22[7] , 
        \R_DATA_TEMPR22[6] , \R_DATA_TEMPR22[5] , \R_DATA_TEMPR22[4] , 
        \R_DATA_TEMPR22[3] , \R_DATA_TEMPR22[2] , \R_DATA_TEMPR22[1] , 
        \R_DATA_TEMPR22[0] }));
    OR4 OR4_245 (.A(OR4_100_Y), .B(OR2_0_Y), .C(\R_DATA_TEMPR22[12] ), 
        .D(\R_DATA_TEMPR23[12] ), .Y(OR4_245_Y));
    OR4 OR4_50 (.A(\R_DATA_TEMPR16[5] ), .B(\R_DATA_TEMPR17[5] ), .C(
        \R_DATA_TEMPR18[5] ), .D(\R_DATA_TEMPR19[5] ), .Y(OR4_50_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R2C3 (.BLK_EN(\BLKX0[2] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][3] ), .R_DATA({nc138, nc139, 
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR2[38] , \R_DATA_TEMPR2[37] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR2[35] , \R_DATA_TEMPR2[34] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR2[32] , \R_DATA_TEMPR2[31] , 
        \R_DATA_TEMPR2[30] }));
    OR4 OR4_57 (.A(\R_DATA_TEMPR0[36] ), .B(\R_DATA_TEMPR1[36] ), .C(
        \R_DATA_TEMPR2[36] ), .D(\R_DATA_TEMPR3[36] ), .Y(OR4_57_Y));
    OR4 OR4_32 (.A(\R_DATA_TEMPR16[20] ), .B(\R_DATA_TEMPR17[20] ), .C(
        \R_DATA_TEMPR18[20] ), .D(\R_DATA_TEMPR19[20] ), .Y(OR4_32_Y));
    OR4 OR4_260 (.A(\R_DATA_TEMPR28[38] ), .B(\R_DATA_TEMPR29[38] ), 
        .C(\R_DATA_TEMPR30[38] ), .D(\R_DATA_TEMPR31[38] ), .Y(
        OR4_260_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[7]  (.A(CFG3_3_Y), .B(CFG3_4_Y), 
        .Y(\BLKZ0[7] ));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R10C3 (.BLK_EN(\BLKX0[10] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][3] ), .R_DATA({nc140, nc141, 
        \R_DATA_TEMPR10[39] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR10[37] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR10[35] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR10[33] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR10[31] , \R_DATA_TEMPR10[30] }));
    OR4 OR4_184 (.A(\R_DATA_TEMPR0[37] ), .B(\R_DATA_TEMPR1[37] ), .C(
        \R_DATA_TEMPR2[37] ), .D(\R_DATA_TEMPR3[37] ), .Y(OR4_184_Y));
    OR4 OR4_311 (.A(OR4_52_Y), .B(OR2_29_Y), .C(\R_DATA_TEMPR22[21] ), 
        .D(\R_DATA_TEMPR23[21] ), .Y(OR4_311_Y));
    OR4 OR4_248 (.A(\R_DATA_TEMPR8[16] ), .B(\R_DATA_TEMPR9[16] ), .C(
        \R_DATA_TEMPR10[16] ), .D(\R_DATA_TEMPR11[16] ), .Y(OR4_248_Y));
    OR4 OR4_302 (.A(\R_DATA_TEMPR4[15] ), .B(\R_DATA_TEMPR5[15] ), .C(
        \R_DATA_TEMPR6[15] ), .D(\R_DATA_TEMPR7[15] ), .Y(OR4_302_Y));
    OR4 OR4_266 (.A(\R_DATA_TEMPR0[10] ), .B(\R_DATA_TEMPR1[10] ), .C(
        \R_DATA_TEMPR2[10] ), .D(\R_DATA_TEMPR3[10] ), .Y(OR4_266_Y));
    OR4 OR4_10 (.A(\R_DATA_TEMPR28[20] ), .B(\R_DATA_TEMPR29[20] ), .C(
        \R_DATA_TEMPR30[20] ), .D(\R_DATA_TEMPR31[20] ), .Y(OR4_10_Y));
    OR4 OR4_25 (.A(\R_DATA_TEMPR16[34] ), .B(\R_DATA_TEMPR17[34] ), .C(
        \R_DATA_TEMPR18[34] ), .D(\R_DATA_TEMPR19[34] ), .Y(OR4_25_Y));
    OR4 OR4_76 (.A(\R_DATA_TEMPR0[27] ), .B(\R_DATA_TEMPR1[27] ), .C(
        \R_DATA_TEMPR2[27] ), .D(\R_DATA_TEMPR3[27] ), .Y(OR4_76_Y));
    OR4 OR4_339 (.A(\R_DATA_TEMPR24[17] ), .B(\R_DATA_TEMPR25[17] ), 
        .C(\R_DATA_TEMPR26[17] ), .D(\R_DATA_TEMPR27[17] ), .Y(
        OR4_339_Y));
    OR4 OR4_193 (.A(OR4_341_Y), .B(OR4_107_Y), .C(OR4_253_Y), .D(
        OR4_38_Y), .Y(OR4_193_Y));
    OR4 OR4_17 (.A(\R_DATA_TEMPR12[34] ), .B(\R_DATA_TEMPR13[34] ), .C(
        \R_DATA_TEMPR14[34] ), .D(\R_DATA_TEMPR15[34] ), .Y(OR4_17_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R24C2 (.BLK_EN(\BLKX0[24] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[24] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][2] ), .R_DATA({nc142, nc143, 
        \R_DATA_TEMPR24[29] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR24[27] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR24[25] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR24[23] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR24[21] , \R_DATA_TEMPR24[20] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R30C0 (.BLK_EN(\BLKX0[30] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[30] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][0] ), .R_DATA({nc144, nc145, 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR30[4] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR30[0] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R2C0 (.BLK_EN(\BLKX0[2] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[2] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][0] ), .R_DATA({nc146, nc147, 
        \R_DATA_TEMPR2[9] , \R_DATA_TEMPR2[8] , \R_DATA_TEMPR2[7] , 
        \R_DATA_TEMPR2[6] , \R_DATA_TEMPR2[5] , \R_DATA_TEMPR2[4] , 
        \R_DATA_TEMPR2[3] , \R_DATA_TEMPR2[2] , \R_DATA_TEMPR2[1] , 
        \R_DATA_TEMPR2[0] }));
    CFG3 #( .INIT(8'h20) )  CFG3_14 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_14_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R31C3 (.BLK_EN(\BLKX0[31] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[31] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][3] ), .R_DATA({nc148, nc149, 
        \R_DATA_TEMPR31[39] , \R_DATA_TEMPR31[38] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR31[36] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR31[34] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR31[32] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR31[30] }));
    OR4 OR4_200 (.A(\R_DATA_TEMPR12[33] ), .B(\R_DATA_TEMPR13[33] ), 
        .C(\R_DATA_TEMPR14[33] ), .D(\R_DATA_TEMPR15[33] ), .Y(
        OR4_200_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R21C1 (.BLK_EN(\BLKX0[21] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[21] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][1] ), .R_DATA({nc150, nc151, 
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR21[18] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR21[16] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR21[14] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR21[12] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR21[10] }));
    OR4 OR4_270 (.A(\R_DATA_TEMPR8[10] ), .B(\R_DATA_TEMPR9[10] ), .C(
        \R_DATA_TEMPR10[10] ), .D(\R_DATA_TEMPR11[10] ), .Y(OR4_270_Y));
    OR4 OR4_319 (.A(\R_DATA_TEMPR8[15] ), .B(\R_DATA_TEMPR9[15] ), .C(
        \R_DATA_TEMPR10[15] ), .D(\R_DATA_TEMPR11[15] ), .Y(OR4_319_Y));
    OR4 OR4_192 (.A(OR4_231_Y), .B(OR4_113_Y), .C(OR4_234_Y), .D(
        OR4_104_Y), .Y(OR4_192_Y));
    OR4 OR4_123 (.A(\R_DATA_TEMPR12[3] ), .B(\R_DATA_TEMPR13[3] ), .C(
        \R_DATA_TEMPR14[3] ), .D(\R_DATA_TEMPR15[3] ), .Y(OR4_123_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R0C1 (.BLK_EN(\BLKX0[0] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][1] ), .R_DATA({nc152, nc153, 
        \R_DATA_TEMPR0[19] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR0[17] , 
        \R_DATA_TEMPR0[16] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR0[14] , 
        \R_DATA_TEMPR0[13] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR0[11] , 
        \R_DATA_TEMPR0[10] }));
    OR4 OR4_206 (.A(OR4_350_Y), .B(OR4_44_Y), .C(OR4_261_Y), .D(
        OR4_215_Y), .Y(OR4_206_Y));
    OR4 OR4_70 (.A(\R_DATA_TEMPR24[31] ), .B(\R_DATA_TEMPR25[31] ), .C(
        \R_DATA_TEMPR26[31] ), .D(\R_DATA_TEMPR27[31] ), .Y(OR4_70_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[17]  (.A(CFG3_0_Y), .B(CFG3_9_Y)
        , .Y(\BLKX0[17] ));
    OR4 OR4_58 (.A(OR4_5_Y), .B(OR4_80_Y), .C(OR4_125_Y), .D(OR4_17_Y), 
        .Y(OR4_58_Y));
    OR4 OR4_276 (.A(\R_DATA_TEMPR4[27] ), .B(\R_DATA_TEMPR5[27] ), .C(
        \R_DATA_TEMPR6[27] ), .D(\R_DATA_TEMPR7[27] ), .Y(OR4_276_Y));
    OR4 OR4_242 (.A(\R_DATA_TEMPR28[35] ), .B(\R_DATA_TEMPR29[35] ), 
        .C(\R_DATA_TEMPR30[35] ), .D(\R_DATA_TEMPR31[35] ), .Y(
        OR4_242_Y));
    OR4 OR4_77 (.A(OR4_109_Y), .B(OR4_303_Y), .C(OR4_81_Y), .D(
        OR4_250_Y), .Y(OR4_77_Y));
    OR4 OR4_299 (.A(OR4_25_Y), .B(OR2_17_Y), .C(\R_DATA_TEMPR22[34] ), 
        .D(\R_DATA_TEMPR23[34] ), .Y(OR4_299_Y));
    OR4 \OR4_R_DATA[5]  (.A(OR4_51_Y), .B(OR4_343_Y), .C(OR4_222_Y), 
        .D(OR4_298_Y), .Y(R_DATA[5]));
    OR4 OR4_340 (.A(\R_DATA_TEMPR0[16] ), .B(\R_DATA_TEMPR1[16] ), .C(
        \R_DATA_TEMPR2[16] ), .D(\R_DATA_TEMPR3[16] ), .Y(OR4_340_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R6C2 (.BLK_EN(\BLKX0[6] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][2] ), .R_DATA({nc154, nc155, 
        \R_DATA_TEMPR6[29] , \R_DATA_TEMPR6[28] , \R_DATA_TEMPR6[27] , 
        \R_DATA_TEMPR6[26] , \R_DATA_TEMPR6[25] , \R_DATA_TEMPR6[24] , 
        \R_DATA_TEMPR6[23] , \R_DATA_TEMPR6[22] , \R_DATA_TEMPR6[21] , 
        \R_DATA_TEMPR6[20] }));
    OR4 \OR4_R_DATA[11]  (.A(OR4_0_Y), .B(OR4_346_Y), .C(OR4_356_Y), 
        .D(OR4_237_Y), .Y(R_DATA[11]));
    OR4 OR4_122 (.A(OR4_277_Y), .B(OR2_32_Y), .C(\R_DATA_TEMPR22[39] ), 
        .D(\R_DATA_TEMPR23[39] ), .Y(OR4_122_Y));
    OR4 \OR4_R_DATA[9]  (.A(OR4_41_Y), .B(OR4_118_Y), .C(OR4_203_Y), 
        .D(OR4_279_Y), .Y(R_DATA[9]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R14C3 (.BLK_EN(\BLKX0[14] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][3] ), .R_DATA({nc156, nc157, 
        \R_DATA_TEMPR14[39] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR14[37] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR14[35] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR14[33] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR14[31] , \R_DATA_TEMPR14[30] }));
    OR4 OR4_18 (.A(\R_DATA_TEMPR4[35] ), .B(\R_DATA_TEMPR5[35] ), .C(
        \R_DATA_TEMPR6[35] ), .D(\R_DATA_TEMPR7[35] ), .Y(OR4_18_Y));
    OR4 OR4_34 (.A(\R_DATA_TEMPR8[35] ), .B(\R_DATA_TEMPR9[35] ), .C(
        \R_DATA_TEMPR10[35] ), .D(\R_DATA_TEMPR11[35] ), .Y(OR4_34_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R22C3 (.BLK_EN(\BLKX0[22] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[22] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][3] ), .R_DATA({nc158, nc159, 
        \R_DATA_TEMPR22[39] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR22[37] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR22[35] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR22[33] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR22[31] , \R_DATA_TEMPR22[30] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R9C3 (.BLK_EN(\BLKX0[9] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][3] ), .R_DATA({nc160, nc161, 
        \R_DATA_TEMPR9[39] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR9[37] , 
        \R_DATA_TEMPR9[36] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR9[34] , 
        \R_DATA_TEMPR9[33] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR9[31] , 
        \R_DATA_TEMPR9[30] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R14C1 (.BLK_EN(\BLKX0[14] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][1] ), .R_DATA({nc162, nc163, 
        \R_DATA_TEMPR14[19] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR14[17] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR14[15] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR14[13] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR14[11] , \R_DATA_TEMPR14[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R8C2 (.BLK_EN(\BLKX0[8] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][2] ), .R_DATA({nc164, nc165, 
        \R_DATA_TEMPR8[29] , \R_DATA_TEMPR8[28] , \R_DATA_TEMPR8[27] , 
        \R_DATA_TEMPR8[26] , \R_DATA_TEMPR8[25] , \R_DATA_TEMPR8[24] , 
        \R_DATA_TEMPR8[23] , \R_DATA_TEMPR8[22] , \R_DATA_TEMPR8[21] , 
        \R_DATA_TEMPR8[20] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R17C2 (.BLK_EN(\BLKX0[17] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][2] ), .R_DATA({nc166, nc167, 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR17[28] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR17[26] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR17[24] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR17[22] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR17[20] }));
    OR4 \OR4_R_DATA[35]  (.A(OR4_27_Y), .B(OR4_204_Y), .C(OR4_352_Y), 
        .D(OR4_242_Y), .Y(R_DATA[35]));
    OR4 \OR4_R_DATA[10]  (.A(OR4_294_Y), .B(OR4_13_Y), .C(OR4_171_Y), 
        .D(OR4_33_Y), .Y(R_DATA[10]));
    OR4 OR4_229 (.A(\R_DATA_TEMPR4[16] ), .B(\R_DATA_TEMPR5[16] ), .C(
        \R_DATA_TEMPR6[16] ), .D(\R_DATA_TEMPR7[16] ), .Y(OR4_229_Y));
    OR4 OR4_356 (.A(\R_DATA_TEMPR24[11] ), .B(\R_DATA_TEMPR25[11] ), 
        .C(\R_DATA_TEMPR26[11] ), .D(\R_DATA_TEMPR27[11] ), .Y(
        OR4_356_Y));
    OR4 OR4_261 (.A(\R_DATA_TEMPR8[7] ), .B(\R_DATA_TEMPR9[7] ), .C(
        \R_DATA_TEMPR10[7] ), .D(\R_DATA_TEMPR11[7] ), .Y(OR4_261_Y));
    OR2 OR2_23 (.A(\R_DATA_TEMPR20[2] ), .B(\R_DATA_TEMPR21[2] ), .Y(
        OR2_23_Y));
    OR4 OR4_29 (.A(\R_DATA_TEMPR28[12] ), .B(\R_DATA_TEMPR29[12] ), .C(
        \R_DATA_TEMPR30[12] ), .D(\R_DATA_TEMPR31[12] ), .Y(OR4_29_Y));
    OR4 \OR4_R_DATA[16]  (.A(OR4_160_Y), .B(OR4_2_Y), .C(OR4_63_Y), .D(
        OR4_86_Y), .Y(R_DATA[16]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R22C2 (.BLK_EN(\BLKX0[22] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[22] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][2] ), .R_DATA({nc168, nc169, 
        \R_DATA_TEMPR22[29] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR22[27] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR22[25] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR22[23] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR22[21] , \R_DATA_TEMPR22[20] }));
    OR4 OR4_280 (.A(\R_DATA_TEMPR28[29] ), .B(\R_DATA_TEMPR29[29] ), 
        .C(\R_DATA_TEMPR30[29] ), .D(\R_DATA_TEMPR31[29] ), .Y(
        OR4_280_Y));
    OR4 OR4_233 (.A(\R_DATA_TEMPR4[23] ), .B(\R_DATA_TEMPR5[23] ), .C(
        \R_DATA_TEMPR6[23] ), .D(\R_DATA_TEMPR7[23] ), .Y(OR4_233_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R22C1 (.BLK_EN(\BLKX0[22] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[22] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][1] ), .R_DATA({nc170, nc171, 
        \R_DATA_TEMPR22[19] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR22[17] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR22[15] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR22[13] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR22[11] , \R_DATA_TEMPR22[10] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[31]  (.A(CFG3_3_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[31] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[25]  (.A(CFG3_0_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[25] ));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R7C1 (.BLK_EN(\BLKX0[7] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][1] ), .R_DATA({nc172, nc173, 
        \R_DATA_TEMPR7[19] , \R_DATA_TEMPR7[18] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR7[16] , \R_DATA_TEMPR7[15] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR7[13] , \R_DATA_TEMPR7[12] , \R_DATA_TEMPR7[11] , 
        \R_DATA_TEMPR7[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R15C1 (.BLK_EN(\BLKX0[15] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][1] ), .R_DATA({nc174, nc175, 
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR15[18] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR15[16] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR15[14] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR15[12] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR15[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R25C2 (.BLK_EN(\BLKX0[25] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[25] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][2] ), .R_DATA({nc176, nc177, 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR25[28] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR25[26] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR25[24] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR25[22] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR25[20] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[20]  (.A(CFG3_18_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[20] ));
    OR4 OR4_286 (.A(\R_DATA_TEMPR0[14] ), .B(\R_DATA_TEMPR1[14] ), .C(
        \R_DATA_TEMPR2[14] ), .D(\R_DATA_TEMPR3[14] ), .Y(OR4_286_Y));
    OR4 OR4_78 (.A(\R_DATA_TEMPR12[9] ), .B(\R_DATA_TEMPR13[9] ), .C(
        \R_DATA_TEMPR14[9] ), .D(\R_DATA_TEMPR15[9] ), .Y(OR4_78_Y));
    OR4 \OR4_R_DATA[8]  (.A(OR4_174_Y), .B(OR4_214_Y), .C(OR4_134_Y), 
        .D(OR4_269_Y), .Y(R_DATA[8]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R20C2 (.BLK_EN(\BLKX0[20] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[20] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][2] ), .R_DATA({nc178, nc179, 
        \R_DATA_TEMPR20[29] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR20[27] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR20[25] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR20[23] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR20[21] , \R_DATA_TEMPR20[20] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R10C0 (.BLK_EN(\BLKX0[10] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][0] ), .R_DATA({nc180, nc181, 
        \R_DATA_TEMPR10[9] , \R_DATA_TEMPR10[8] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR10[6] , \R_DATA_TEMPR10[5] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR10[3] , \R_DATA_TEMPR10[2] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR10[0] }));
    OR4 OR4_154 (.A(\R_DATA_TEMPR4[20] ), .B(\R_DATA_TEMPR5[20] ), .C(
        \R_DATA_TEMPR6[20] ), .D(\R_DATA_TEMPR7[20] ), .Y(OR4_154_Y));
    OR2 OR2_21 (.A(\R_DATA_TEMPR20[8] ), .B(\R_DATA_TEMPR21[8] ), .Y(
        OR2_21_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R11C3 (.BLK_EN(\BLKX0[11] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][3] ), .R_DATA({nc182, nc183, 
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR11[38] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR11[36] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR11[34] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR11[32] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR11[30] }));
    OR4 OR4_22 (.A(\R_DATA_TEMPR28[39] ), .B(\R_DATA_TEMPR29[39] ), .C(
        \R_DATA_TEMPR30[39] ), .D(\R_DATA_TEMPR31[39] ), .Y(OR4_22_Y));
    OR4 OR4_143 (.A(\R_DATA_TEMPR28[28] ), .B(\R_DATA_TEMPR29[28] ), 
        .C(\R_DATA_TEMPR30[28] ), .D(\R_DATA_TEMPR31[28] ), .Y(
        OR4_143_Y));
    OR4 OR4_213 (.A(OR4_62_Y), .B(OR2_16_Y), .C(\R_DATA_TEMPR22[22] ), 
        .D(\R_DATA_TEMPR23[22] ), .Y(OR4_213_Y));
    OR4 OR4_201 (.A(\R_DATA_TEMPR0[31] ), .B(\R_DATA_TEMPR1[31] ), .C(
        \R_DATA_TEMPR2[31] ), .D(\R_DATA_TEMPR3[31] ), .Y(OR4_201_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R16C3 (.BLK_EN(\BLKX0[16] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][3] ), .R_DATA({nc184, nc185, 
        \R_DATA_TEMPR16[39] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR16[37] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR16[35] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR16[33] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR16[31] , \R_DATA_TEMPR16[30] }));
    OR2 OR2_13 (.A(\R_DATA_TEMPR20[18] ), .B(\R_DATA_TEMPR21[18] ), .Y(
        OR2_13_Y));
    OR4 OR4_6 (.A(\R_DATA_TEMPR12[1] ), .B(\R_DATA_TEMPR13[1] ), .C(
        \R_DATA_TEMPR14[1] ), .D(\R_DATA_TEMPR15[1] ), .Y(OR4_6_Y));
    OR4 OR4_271 (.A(\R_DATA_TEMPR28[34] ), .B(\R_DATA_TEMPR29[34] ), 
        .C(\R_DATA_TEMPR30[34] ), .D(\R_DATA_TEMPR31[34] ), .Y(
        OR4_271_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R13C2 (.BLK_EN(\BLKX0[13] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][2] ), .R_DATA({nc186, nc187, 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR13[28] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR13[26] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR13[24] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR13[22] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR13[20] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[3]  (.A(CFG3_19_Y), .B(CFG3_5_Y)
        , .Y(\BLKX0[3] ));
    CFG3 #( .INIT(8'h4) )  CFG3_8 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_8_Y));
    OR4 \OR4_R_DATA[17]  (.A(OR4_77_Y), .B(OR4_244_Y), .C(OR4_339_Y), 
        .D(OR4_12_Y), .Y(R_DATA[17]));
    OR4 OR4_142 (.A(\R_DATA_TEMPR24[36] ), .B(\R_DATA_TEMPR25[36] ), 
        .C(\R_DATA_TEMPR26[36] ), .D(\R_DATA_TEMPR27[36] ), .Y(
        OR4_142_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[23]  (.A(CFG3_3_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[23] ));
    OR2 OR2_11 (.A(\R_DATA_TEMPR20[30] ), .B(\R_DATA_TEMPR21[30] ), .Y(
        OR2_11_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[2]  (.A(CFG3_8_Y), .B(CFG3_5_Y), 
        .Y(\BLKX0[2] ));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R31C1 (.BLK_EN(\BLKX0[31] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[31] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][1] ), .R_DATA({nc188, nc189, 
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR31[18] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR31[16] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR31[14] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR31[12] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR31[10] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R28C3 (.BLK_EN(\BLKX0[28] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[28] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][3] ), .R_DATA({nc190, nc191, 
        \R_DATA_TEMPR28[39] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR28[37] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR28[35] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR28[33] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR28[31] , \R_DATA_TEMPR28[30] }));
    OR4 OR4_55 (.A(\R_DATA_TEMPR28[6] ), .B(\R_DATA_TEMPR29[6] ), .C(
        \R_DATA_TEMPR30[6] ), .D(\R_DATA_TEMPR31[6] ), .Y(OR4_55_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[5]  (.A(CFG3_14_Y), .B(CFG3_4_Y)
        , .Y(\BLKZ0[5] ));
    OR4 OR4_301 (.A(OR4_54_Y), .B(OR4_357_Y), .C(OR4_348_Y), .D(
        OR4_200_Y), .Y(OR4_301_Y));
    OR4 OR4_249 (.A(\R_DATA_TEMPR0[24] ), .B(\R_DATA_TEMPR1[24] ), .C(
        \R_DATA_TEMPR2[24] ), .D(\R_DATA_TEMPR3[24] ), .Y(OR4_249_Y));
    OR4 \OR4_R_DATA[38]  (.A(OR4_60_Y), .B(OR4_15_Y), .C(OR4_208_Y), 
        .D(OR4_260_Y), .Y(R_DATA[38]));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[19]  (.A(CFG3_19_Y), .B(
        CFG3_9_Y), .Y(\BLKX0[19] ));
    OR4 OR4_352 (.A(\R_DATA_TEMPR24[35] ), .B(\R_DATA_TEMPR25[35] ), 
        .C(\R_DATA_TEMPR26[35] ), .D(\R_DATA_TEMPR27[35] ), .Y(
        OR4_352_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[15]  (.A(CFG3_3_Y), .B(
        CFG3_20_Y), .Y(\BLKZ0[15] ));
    OR4 OR4_15 (.A(OR4_183_Y), .B(OR2_18_Y), .C(\R_DATA_TEMPR22[38] ), 
        .D(\R_DATA_TEMPR23[38] ), .Y(OR4_15_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R15C3 (.BLK_EN(\BLKX0[15] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][3] ), .R_DATA({nc192, nc193, 
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR15[38] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR15[36] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR15[34] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR15[32] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR15[30] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R24C0 (.BLK_EN(\BLKX0[24] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[24] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][0] ), .R_DATA({nc194, nc195, 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR24[4] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR24[1] , 
        \R_DATA_TEMPR24[0] }));
    OR4 OR4_281 (.A(\R_DATA_TEMPR16[37] ), .B(\R_DATA_TEMPR17[37] ), 
        .C(\R_DATA_TEMPR18[37] ), .D(\R_DATA_TEMPR19[37] ), .Y(
        OR4_281_Y));
    OR4 OR4_326 (.A(\R_DATA_TEMPR0[1] ), .B(\R_DATA_TEMPR1[1] ), .C(
        \R_DATA_TEMPR2[1] ), .D(\R_DATA_TEMPR3[1] ), .Y(OR4_326_Y));
    OR4 OR4_194 (.A(\R_DATA_TEMPR12[38] ), .B(\R_DATA_TEMPR13[38] ), 
        .C(\R_DATA_TEMPR14[38] ), .D(\R_DATA_TEMPR15[38] ), .Y(
        OR4_194_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R5C0 (.BLK_EN(\BLKX0[5] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][0] ), .R_DATA({nc196, nc197, 
        \R_DATA_TEMPR5[9] , \R_DATA_TEMPR5[8] , \R_DATA_TEMPR5[7] , 
        \R_DATA_TEMPR5[6] , \R_DATA_TEMPR5[5] , \R_DATA_TEMPR5[4] , 
        \R_DATA_TEMPR5[3] , \R_DATA_TEMPR5[2] , \R_DATA_TEMPR5[1] , 
        \R_DATA_TEMPR5[0] }));
    OR4 OR4_93 (.A(\R_DATA_TEMPR12[23] ), .B(\R_DATA_TEMPR13[23] ), .C(
        \R_DATA_TEMPR14[23] ), .D(\R_DATA_TEMPR15[23] ), .Y(OR4_93_Y));
    OR4 OR4_309 (.A(\R_DATA_TEMPR16[14] ), .B(\R_DATA_TEMPR17[14] ), 
        .C(\R_DATA_TEMPR18[14] ), .D(\R_DATA_TEMPR19[14] ), .Y(
        OR4_309_Y));
    OR4 OR4_24 (.A(\R_DATA_TEMPR8[1] ), .B(\R_DATA_TEMPR9[1] ), .C(
        \R_DATA_TEMPR10[1] ), .D(\R_DATA_TEMPR11[1] ), .Y(OR4_24_Y));
    OR4 OR4_8 (.A(\R_DATA_TEMPR8[24] ), .B(\R_DATA_TEMPR9[24] ), .C(
        \R_DATA_TEMPR10[24] ), .D(\R_DATA_TEMPR11[24] ), .Y(OR4_8_Y));
    OR4 OR4_250 (.A(\R_DATA_TEMPR12[17] ), .B(\R_DATA_TEMPR13[17] ), 
        .C(\R_DATA_TEMPR14[17] ), .D(\R_DATA_TEMPR15[17] ), .Y(
        OR4_250_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R13C1 (.BLK_EN(\BLKX0[13] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][1] ), .R_DATA({nc198, nc199, 
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR13[18] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR13[16] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR13[14] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR13[12] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR13[10] }));
    OR4 OR4_334 (.A(OR4_209_Y), .B(OR2_34_Y), .C(\R_DATA_TEMPR22[1] ), 
        .D(\R_DATA_TEMPR23[1] ), .Y(OR4_334_Y));
    OR2 OR2_4 (.A(\R_DATA_TEMPR20[10] ), .B(\R_DATA_TEMPR21[10] ), .Y(
        OR2_4_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R17C0 (.BLK_EN(\BLKX0[17] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][0] ), .R_DATA({nc200, nc201, 
        \R_DATA_TEMPR17[9] , \R_DATA_TEMPR17[8] , \R_DATA_TEMPR17[7] , 
        \R_DATA_TEMPR17[6] , \R_DATA_TEMPR17[5] , \R_DATA_TEMPR17[4] , 
        \R_DATA_TEMPR17[3] , \R_DATA_TEMPR17[2] , \R_DATA_TEMPR17[1] , 
        \R_DATA_TEMPR17[0] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R12C0 (.BLK_EN(\BLKX0[12] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][0] ), .R_DATA({nc202, nc203, 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR12[0] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R27C1 (.BLK_EN(\BLKX0[27] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[27] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][1] ), .R_DATA({nc204, nc205, 
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR27[18] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR27[16] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR27[14] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR27[12] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR27[10] }));
    OR4 OR4_131 (.A(\R_DATA_TEMPR4[28] ), .B(\R_DATA_TEMPR5[28] ), .C(
        \R_DATA_TEMPR6[28] ), .D(\R_DATA_TEMPR7[28] ), .Y(OR4_131_Y));
    OR4 \OR4_R_DATA[39]  (.A(OR4_193_Y), .B(OR4_122_Y), .C(OR4_95_Y), 
        .D(OR4_22_Y), .Y(R_DATA[39]));
    OR4 OR4_256 (.A(OR4_324_Y), .B(OR4_169_Y), .C(OR4_247_Y), .D(
        OR4_72_Y), .Y(OR4_256_Y));
    OR2 OR2_0 (.A(\R_DATA_TEMPR20[12] ), .B(\R_DATA_TEMPR21[12] ), .Y(
        OR2_0_Y));
    OR4 OR4_75 (.A(\R_DATA_TEMPR4[8] ), .B(\R_DATA_TEMPR5[8] ), .C(
        \R_DATA_TEMPR6[8] ), .D(\R_DATA_TEMPR7[8] ), .Y(OR4_75_Y));
    OR2 OR2_6 (.A(\R_DATA_TEMPR20[32] ), .B(\R_DATA_TEMPR21[32] ), .Y(
        OR2_6_Y));
    OR4 OR4_91 (.A(\R_DATA_TEMPR16[16] ), .B(\R_DATA_TEMPR17[16] ), .C(
        \R_DATA_TEMPR18[16] ), .D(\R_DATA_TEMPR19[16] ), .Y(OR4_91_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_2 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_2_Y));
    OR4 OR4_124 (.A(\R_DATA_TEMPR28[32] ), .B(\R_DATA_TEMPR29[32] ), 
        .C(\R_DATA_TEMPR30[32] ), .D(\R_DATA_TEMPR31[32] ), .Y(
        OR4_124_Y));
    OR2 OR2_3 (.A(\R_DATA_TEMPR20[9] ), .B(\R_DATA_TEMPR21[9] ), .Y(
        OR2_3_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R21C2 (.BLK_EN(\BLKX0[21] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[21] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][2] ), .R_DATA({nc206, nc207, 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR21[28] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR21[26] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR21[24] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR21[22] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR21[20] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[4]  (.A(CFG3_21_Y), .B(CFG3_5_Y)
        , .Y(\BLKX0[4] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[21]  (.A(CFG3_14_Y), .B(
        CFG3_13_Y), .Y(\BLKZ0[21] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[26]  (.A(CFG3_16_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[26] ));
    OR4 OR4_314 (.A(\R_DATA_TEMPR0[38] ), .B(\R_DATA_TEMPR1[38] ), .C(
        \R_DATA_TEMPR2[38] ), .D(\R_DATA_TEMPR3[38] ), .Y(OR4_314_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_21 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_21_Y));
    OR4 OR4_43 (.A(\R_DATA_TEMPR0[6] ), .B(\R_DATA_TEMPR1[6] ), .C(
        \R_DATA_TEMPR2[6] ), .D(\R_DATA_TEMPR3[6] ), .Y(OR4_43_Y));
    OR2 OR2_26 (.A(\R_DATA_TEMPR20[24] ), .B(\R_DATA_TEMPR21[24] ), .Y(
        OR2_26_Y));
    OR4 OR4_111 (.A(\R_DATA_TEMPR4[4] ), .B(\R_DATA_TEMPR5[4] ), .C(
        \R_DATA_TEMPR6[4] ), .D(\R_DATA_TEMPR7[4] ), .Y(OR4_111_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_1 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_1_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R5C3 (.BLK_EN(\BLKX0[5] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][3] ), .R_DATA({nc208, nc209, 
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR5[38] , \R_DATA_TEMPR5[37] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR5[35] , \R_DATA_TEMPR5[34] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR5[32] , \R_DATA_TEMPR5[31] , 
        \R_DATA_TEMPR5[30] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R30C2 (.BLK_EN(\BLKX0[30] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[30] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][2] ), .R_DATA({nc210, nc211, 
        \R_DATA_TEMPR30[29] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR30[27] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR30[25] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR30[23] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR30[21] , \R_DATA_TEMPR30[20] }));
    OR4 OR4_59 (.A(\R_DATA_TEMPR0[25] ), .B(\R_DATA_TEMPR1[25] ), .C(
        \R_DATA_TEMPR2[25] ), .D(\R_DATA_TEMPR3[25] ), .Y(OR4_59_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R14C2 (.BLK_EN(\BLKX0[14] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][2] ), .R_DATA({nc212, nc213, 
        \R_DATA_TEMPR14[29] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR14[27] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR14[25] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR14[23] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR14[21] , \R_DATA_TEMPR14[20] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R1C0 (.BLK_EN(\BLKX0[1] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][0] ), .R_DATA({nc214, nc215, 
        \R_DATA_TEMPR1[9] , \R_DATA_TEMPR1[8] , \R_DATA_TEMPR1[7] , 
        \R_DATA_TEMPR1[6] , \R_DATA_TEMPR1[5] , \R_DATA_TEMPR1[4] , 
        \R_DATA_TEMPR1[3] , \R_DATA_TEMPR1[2] , \R_DATA_TEMPR1[1] , 
        \R_DATA_TEMPR1[0] }));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R8C1 (.BLK_EN(\BLKX0[8] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][1] ), .R_DATA({nc216, nc217, 
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR8[18] , \R_DATA_TEMPR8[17] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR8[15] , \R_DATA_TEMPR8[14] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR8[12] , \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR8[10] }));
    OR4 OR4_263 (.A(\R_DATA_TEMPR24[15] ), .B(\R_DATA_TEMPR25[15] ), 
        .C(\R_DATA_TEMPR26[15] ), .D(\R_DATA_TEMPR27[15] ), .Y(
        OR4_263_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[14]  (.A(CFG3_7_Y), .B(
        CFG3_20_Y), .Y(\BLKZ0[14] ));
    CFG3 #( .INIT(8'h1) )  CFG3_11 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_11_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R28C2 (.BLK_EN(\BLKX0[28] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[28] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][2] ), .R_DATA({nc218, nc219, 
        \R_DATA_TEMPR28[29] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR28[27] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR28[25] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR28[23] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR28[21] , \R_DATA_TEMPR28[20] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[22]  (.A(CFG3_2_Y), .B(CFG3_9_Y)
        , .Y(\BLKX0[22] ));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R11C1 (.BLK_EN(\BLKX0[11] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][1] ), .R_DATA({nc220, nc221, 
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR11[18] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR11[16] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR11[14] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR11[12] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR11[10] }));
    OR4 \OR4_R_DATA[0]  (.A(OR4_297_Y), .B(OR4_337_Y), .C(OR4_220_Y), 
        .D(OR4_293_Y), .Y(R_DATA[0]));
    OR4 OR4_19 (.A(\R_DATA_TEMPR4[37] ), .B(\R_DATA_TEMPR5[37] ), .C(
        \R_DATA_TEMPR6[37] ), .D(\R_DATA_TEMPR7[37] ), .Y(OR4_19_Y));
    OR4 OR4_333 (.A(\R_DATA_TEMPR8[36] ), .B(\R_DATA_TEMPR9[36] ), .C(
        \R_DATA_TEMPR10[36] ), .D(\R_DATA_TEMPR11[36] ), .Y(OR4_333_Y));
    OR4 OR4_41 (.A(OR4_116_Y), .B(OR4_315_Y), .C(OR4_197_Y), .D(
        OR4_78_Y), .Y(OR4_41_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[11]  (.A(CFG3_19_Y), .B(
        CFG3_17_Y), .Y(\BLKX0[11] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[30]  (.A(CFG3_2_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[30] ));
    OR4 OR4_52 (.A(\R_DATA_TEMPR16[21] ), .B(\R_DATA_TEMPR17[21] ), .C(
        \R_DATA_TEMPR18[21] ), .D(\R_DATA_TEMPR19[21] ), .Y(OR4_52_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R8C3 (.BLK_EN(\BLKX0[8] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][3] ), .R_DATA({nc222, nc223, 
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR8[38] , \R_DATA_TEMPR8[37] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR8[35] , \R_DATA_TEMPR8[34] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR8[32] , \R_DATA_TEMPR8[31] , 
        \R_DATA_TEMPR8[30] }));
    CFG3 #( .INIT(8'h2) )  CFG3_18 (.A(W_ADDR[8]), .B(W_ADDR[7]), .C(
        W_ADDR[6]), .Y(CFG3_18_Y));
    OR4 OR4_346 (.A(OR4_92_Y), .B(OR2_15_Y), .C(\R_DATA_TEMPR22[11] ), 
        .D(\R_DATA_TEMPR23[11] ), .Y(OR4_346_Y));
    OR4 OR4_136 (.A(\R_DATA_TEMPR12[15] ), .B(\R_DATA_TEMPR13[15] ), 
        .C(\R_DATA_TEMPR14[15] ), .D(\R_DATA_TEMPR15[15] ), .Y(
        OR4_136_Y));
    OR2 OR2_20 (.A(\R_DATA_TEMPR20[20] ), .B(\R_DATA_TEMPR21[20] ), .Y(
        OR2_20_Y));
    OR2 OR2_16 (.A(\R_DATA_TEMPR20[22] ), .B(\R_DATA_TEMPR21[22] ), .Y(
        OR2_16_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_22 (.A(BLK_EN), .B(R_ADDR[10]), .C(
        R_ADDR[9]), .Y(CFG3_22_Y));
    OR2 OR2_27 (.A(\R_DATA_TEMPR20[28] ), .B(\R_DATA_TEMPR21[28] ), .Y(
        OR2_27_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R7C2 (.BLK_EN(\BLKX0[7] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][2] ), .R_DATA({nc224, nc225, 
        \R_DATA_TEMPR7[29] , \R_DATA_TEMPR7[28] , \R_DATA_TEMPR7[27] , 
        \R_DATA_TEMPR7[26] , \R_DATA_TEMPR7[25] , \R_DATA_TEMPR7[24] , 
        \R_DATA_TEMPR7[23] , \R_DATA_TEMPR7[22] , \R_DATA_TEMPR7[21] , 
        \R_DATA_TEMPR7[20] }));
    OR4 OR4_203 (.A(\R_DATA_TEMPR24[9] ), .B(\R_DATA_TEMPR25[9] ), .C(
        \R_DATA_TEMPR26[9] ), .D(\R_DATA_TEMPR27[9] ), .Y(OR4_203_Y));
    OR4 OR4_290 (.A(\R_DATA_TEMPR8[25] ), .B(\R_DATA_TEMPR9[25] ), .C(
        \R_DATA_TEMPR10[25] ), .D(\R_DATA_TEMPR11[25] ), .Y(OR4_290_Y));
    OR4 OR4_338 (.A(\R_DATA_TEMPR24[29] ), .B(\R_DATA_TEMPR25[29] ), 
        .C(\R_DATA_TEMPR26[29] ), .D(\R_DATA_TEMPR27[29] ), .Y(
        OR4_338_Y));
    OR4 OR4_273 (.A(\R_DATA_TEMPR12[24] ), .B(\R_DATA_TEMPR13[24] ), 
        .C(\R_DATA_TEMPR14[24] ), .D(\R_DATA_TEMPR15[24] ), .Y(
        OR4_273_Y));
    OR4 OR4_322 (.A(\R_DATA_TEMPR12[19] ), .B(\R_DATA_TEMPR13[19] ), 
        .C(\R_DATA_TEMPR14[19] ), .D(\R_DATA_TEMPR15[19] ), .Y(
        OR4_322_Y));
    OR4 OR4_313 (.A(\R_DATA_TEMPR16[25] ), .B(\R_DATA_TEMPR17[25] ), 
        .C(\R_DATA_TEMPR18[25] ), .D(\R_DATA_TEMPR19[25] ), .Y(
        OR4_313_Y));
    OR4 OR4_12 (.A(\R_DATA_TEMPR28[17] ), .B(\R_DATA_TEMPR29[17] ), .C(
        \R_DATA_TEMPR30[17] ), .D(\R_DATA_TEMPR31[17] ), .Y(OR4_12_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_12 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_12_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R12C3 (.BLK_EN(\BLKX0[12] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][3] ), .R_DATA({nc226, nc227, 
        \R_DATA_TEMPR12[39] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR12[37] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR12[35] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR12[33] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR12[31] , \R_DATA_TEMPR12[30] }));
    OR4 OR4_296 (.A(\R_DATA_TEMPR0[22] ), .B(\R_DATA_TEMPR1[22] ), .C(
        \R_DATA_TEMPR2[22] ), .D(\R_DATA_TEMPR3[22] ), .Y(OR4_296_Y));
    OR4 OR4_251 (.A(OR4_69_Y), .B(OR2_8_Y), .C(\R_DATA_TEMPR22[6] ), 
        .D(\R_DATA_TEMPR23[6] ), .Y(OR4_251_Y));
    OR4 OR4_79 (.A(\R_DATA_TEMPR24[23] ), .B(\R_DATA_TEMPR25[23] ), .C(
        \R_DATA_TEMPR26[23] ), .D(\R_DATA_TEMPR27[23] ), .Y(OR4_79_Y));
    CFG3 #( .INIT(8'h40) )  CFG3_19 (.A(R_ADDR[8]), .B(R_ADDR[7]), .C(
        R_ADDR[6]), .Y(CFG3_19_Y));
    OR4 OR4_139 (.A(\R_DATA_TEMPR16[3] ), .B(\R_DATA_TEMPR17[3] ), .C(
        \R_DATA_TEMPR18[3] ), .D(\R_DATA_TEMPR19[3] ), .Y(OR4_139_Y));
    OR4 OR4_116 (.A(\R_DATA_TEMPR0[9] ), .B(\R_DATA_TEMPR1[9] ), .C(
        \R_DATA_TEMPR2[9] ), .D(\R_DATA_TEMPR3[9] ), .Y(OR4_116_Y));
    OR4 OR4_144 (.A(\R_DATA_TEMPR16[30] ), .B(\R_DATA_TEMPR17[30] ), 
        .C(\R_DATA_TEMPR18[30] ), .D(\R_DATA_TEMPR19[30] ), .Y(
        OR4_144_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R6C0 (.BLK_EN(\BLKX0[6] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[6] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][0] ), .R_DATA({nc228, nc229, 
        \R_DATA_TEMPR6[9] , \R_DATA_TEMPR6[8] , \R_DATA_TEMPR6[7] , 
        \R_DATA_TEMPR6[6] , \R_DATA_TEMPR6[5] , \R_DATA_TEMPR6[4] , 
        \R_DATA_TEMPR6[3] , \R_DATA_TEMPR6[2] , \R_DATA_TEMPR6[1] , 
        \R_DATA_TEMPR6[0] }));
    OR4 \OR4_R_DATA[32]  (.A(OR4_345_Y), .B(OR4_330_Y), .C(OR4_282_Y), 
        .D(OR4_124_Y), .Y(R_DATA[32]));
    OR4 OR4_220 (.A(\R_DATA_TEMPR24[0] ), .B(\R_DATA_TEMPR25[0] ), .C(
        \R_DATA_TEMPR26[0] ), .D(\R_DATA_TEMPR27[0] ), .Y(OR4_220_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R12C2 (.BLK_EN(\BLKX0[12] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][2] ), .R_DATA({nc230, nc231, 
        \R_DATA_TEMPR12[29] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR12[27] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR12[25] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR12[23] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR12[21] , \R_DATA_TEMPR12[20] }));
    OR4 OR4_318 (.A(\R_DATA_TEMPR12[16] ), .B(\R_DATA_TEMPR13[16] ), 
        .C(\R_DATA_TEMPR14[16] ), .D(\R_DATA_TEMPR15[16] ), .Y(
        OR4_318_Y));
    OR2 OR2_10 (.A(\R_DATA_TEMPR20[23] ), .B(\R_DATA_TEMPR21[23] ), .Y(
        OR2_10_Y));
    OR4 \OR4_R_DATA[3]  (.A(OR4_89_Y), .B(OR4_180_Y), .C(OR4_151_Y), 
        .D(OR4_179_Y), .Y(R_DATA[3]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R12C1 (.BLK_EN(\BLKX0[12] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][1] ), .R_DATA({nc232, nc233, 
        \R_DATA_TEMPR12[19] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR12[17] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR12[15] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR12[13] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR12[11] , \R_DATA_TEMPR12[10] }));
    OR2 OR2_17 (.A(\R_DATA_TEMPR20[34] ), .B(\R_DATA_TEMPR21[34] ), .Y(
        OR2_17_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R15C2 (.BLK_EN(\BLKX0[15] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][2] ), .R_DATA({nc234, nc235, 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR15[28] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR15[26] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR15[24] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR15[22] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR15[20] }));
    OR4 OR4_226 (.A(\R_DATA_TEMPR12[4] ), .B(\R_DATA_TEMPR13[4] ), .C(
        \R_DATA_TEMPR14[4] ), .D(\R_DATA_TEMPR15[4] ), .Y(OR4_226_Y));
    OR4 OR4_119 (.A(\R_DATA_TEMPR24[34] ), .B(\R_DATA_TEMPR25[34] ), 
        .C(\R_DATA_TEMPR26[34] ), .D(\R_DATA_TEMPR27[34] ), .Y(
        OR4_119_Y));
    OR4 OR4_72 (.A(\R_DATA_TEMPR12[12] ), .B(\R_DATA_TEMPR13[12] ), .C(
        \R_DATA_TEMPR14[12] ), .D(\R_DATA_TEMPR15[12] ), .Y(OR4_72_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[24]  (.A(CFG3_6_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[24] ));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R10C2 (.BLK_EN(\BLKX0[10] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][2] ), .R_DATA({nc236, nc237, 
        \R_DATA_TEMPR10[29] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR10[27] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR10[25] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR10[23] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR10[21] , \R_DATA_TEMPR10[20] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[28]  (.A(CFG3_18_Y), .B(
        CFG3_10_Y), .Y(\BLKZ0[28] ));
    OR4 OR4_351 (.A(OR4_32_Y), .B(OR2_20_Y), .C(\R_DATA_TEMPR22[20] ), 
        .D(\R_DATA_TEMPR23[20] ), .Y(OR4_351_Y));
    OR2 OR2_28 (.A(\R_DATA_TEMPR20[19] ), .B(\R_DATA_TEMPR21[19] ), .Y(
        OR2_28_Y));
    OR4 \OR4_R_DATA[33]  (.A(OR4_301_Y), .B(OR4_205_Y), .C(OR4_191_Y), 
        .D(OR4_176_Y), .Y(R_DATA[33]));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R9C1 (.BLK_EN(\BLKX0[9] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][1] ), .R_DATA({nc238, nc239, 
        \R_DATA_TEMPR9[19] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR9[17] , 
        \R_DATA_TEMPR9[16] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR9[14] , 
        \R_DATA_TEMPR9[13] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR9[11] , 
        \R_DATA_TEMPR9[10] }));
    OR4 \OR4_R_DATA[25]  (.A(OR4_285_Y), .B(OR4_97_Y), .C(OR4_230_Y), 
        .D(OR4_133_Y), .Y(R_DATA[25]));
    OR4 OR4_283 (.A(\R_DATA_TEMPR4[0] ), .B(\R_DATA_TEMPR5[0] ), .C(
        \R_DATA_TEMPR6[0] ), .D(\R_DATA_TEMPR7[0] ), .Y(OR4_283_Y));
    OR4 OR4_96 (.A(\R_DATA_TEMPR0[15] ), .B(\R_DATA_TEMPR1[15] ), .C(
        \R_DATA_TEMPR2[15] ), .D(\R_DATA_TEMPR3[15] ), .Y(OR4_96_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_17 (.A(BLK_EN), .B(R_ADDR[10]), .C(
        R_ADDR[9]), .Y(CFG3_17_Y));
    OR4 OR4_54 (.A(\R_DATA_TEMPR0[33] ), .B(\R_DATA_TEMPR1[33] ), .C(
        \R_DATA_TEMPR2[33] ), .D(\R_DATA_TEMPR3[33] ), .Y(OR4_54_Y));
    OR4 OR4_3 (.A(OR4_155_Y), .B(OR2_39_Y), .C(\R_DATA_TEMPR22[29] ), 
        .D(\R_DATA_TEMPR23[29] ), .Y(OR4_3_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R31C2 (.BLK_EN(\BLKX0[31] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[31] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][2] ), .R_DATA({nc240, nc241, 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR31[28] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR31[26] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR31[24] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR31[22] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR31[20] }));
    OR4 OR4_161 (.A(\R_DATA_TEMPR16[27] ), .B(\R_DATA_TEMPR17[27] ), 
        .C(\R_DATA_TEMPR18[27] ), .D(\R_DATA_TEMPR19[27] ), .Y(
        OR4_161_Y));
    OR4 OR4_237 (.A(\R_DATA_TEMPR28[11] ), .B(\R_DATA_TEMPR29[11] ), 
        .C(\R_DATA_TEMPR30[11] ), .D(\R_DATA_TEMPR31[11] ), .Y(
        OR4_237_Y));
    OR4 OR4_137 (.A(\R_DATA_TEMPR16[33] ), .B(\R_DATA_TEMPR17[33] ), 
        .C(\R_DATA_TEMPR18[33] ), .D(\R_DATA_TEMPR19[33] ), .Y(
        OR4_137_Y));
    OR4 OR4_342 (.A(OR4_286_Y), .B(OR4_359_Y), .C(OR4_30_Y), .D(
        OR4_300_Y), .Y(OR4_342_Y));
    OR4 OR4_359 (.A(\R_DATA_TEMPR4[14] ), .B(\R_DATA_TEMPR5[14] ), .C(
        \R_DATA_TEMPR6[14] ), .D(\R_DATA_TEMPR7[14] ), .Y(OR4_359_Y));
    OR4 OR4_14 (.A(OR4_354_Y), .B(OR4_272_Y), .C(OR4_358_Y), .D(
        OR4_148_Y), .Y(OR4_14_Y));
    OR2 OR2_18 (.A(\R_DATA_TEMPR20[38] ), .B(\R_DATA_TEMPR21[38] ), .Y(
        OR2_18_Y));
    OR4 OR4_291 (.A(\R_DATA_TEMPR12[29] ), .B(\R_DATA_TEMPR13[29] ), 
        .C(\R_DATA_TEMPR14[29] ), .D(\R_DATA_TEMPR15[29] ), .Y(
        OR4_291_Y));
    OR4 OR4_234 (.A(\R_DATA_TEMPR8[2] ), .B(\R_DATA_TEMPR9[2] ), .C(
        \R_DATA_TEMPR10[2] ), .D(\R_DATA_TEMPR11[2] ), .Y(OR4_234_Y));
    OR4 OR4_90 (.A(\R_DATA_TEMPR8[6] ), .B(\R_DATA_TEMPR9[6] ), .C(
        \R_DATA_TEMPR10[6] ), .D(\R_DATA_TEMPR11[6] ), .Y(OR4_90_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R18C3 (.BLK_EN(\BLKX0[18] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[39], W_DATA[38], 
        W_DATA[37], W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], 
        W_DATA[32], W_DATA[31], W_DATA[30]}), .W_EN(\BLKZ0[18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][3] ), .R_DATA({nc242, nc243, 
        \R_DATA_TEMPR18[39] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR18[37] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR18[35] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR18[33] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR18[31] , \R_DATA_TEMPR18[30] }));
    OR4 OR4_46 (.A(\R_DATA_TEMPR16[0] ), .B(\R_DATA_TEMPR17[0] ), .C(
        \R_DATA_TEMPR18[0] ), .D(\R_DATA_TEMPR19[0] ), .Y(OR4_46_Y));
    OR4 OR4_97 (.A(OR4_313_Y), .B(OR2_22_Y), .C(\R_DATA_TEMPR22[25] ), 
        .D(\R_DATA_TEMPR23[25] ), .Y(OR4_97_Y));
    OR4 \OR4_R_DATA[6]  (.A(OR4_82_Y), .B(OR4_251_Y), .C(OR4_11_Y), .D(
        OR4_55_Y), .Y(R_DATA[6]));
    OR4 OR4_63 (.A(\R_DATA_TEMPR24[16] ), .B(\R_DATA_TEMPR25[16] ), .C(
        \R_DATA_TEMPR26[16] ), .D(\R_DATA_TEMPR27[16] ), .Y(OR4_63_Y));
    OR4 OR4_217 (.A(\R_DATA_TEMPR8[26] ), .B(\R_DATA_TEMPR9[26] ), .C(
        \R_DATA_TEMPR10[26] ), .D(\R_DATA_TEMPR11[26] ), .Y(OR4_217_Y));
    OR4 OR4_240 (.A(\R_DATA_TEMPR16[2] ), .B(\R_DATA_TEMPR17[2] ), .C(
        \R_DATA_TEMPR18[2] ), .D(\R_DATA_TEMPR19[2] ), .Y(OR4_240_Y));
    OR4 OR4_304 (.A(\R_DATA_TEMPR28[19] ), .B(\R_DATA_TEMPR29[19] ), 
        .C(\R_DATA_TEMPR30[19] ), .D(\R_DATA_TEMPR31[19] ), .Y(
        OR4_304_Y));
    OR4 OR4_117 (.A(OR4_254_Y), .B(OR4_16_Y), .C(OR4_166_Y), .D(
        OR4_322_Y), .Y(OR4_117_Y));
    OR4 OR4_335 (.A(\R_DATA_TEMPR12[37] ), .B(\R_DATA_TEMPR13[37] ), 
        .C(\R_DATA_TEMPR14[37] ), .D(\R_DATA_TEMPR15[37] ), .Y(
        OR4_335_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[20]  (.A(CFG3_21_Y), .B(
        CFG3_9_Y), .Y(\BLKX0[20] ));
    OR4 \OR4_R_DATA[1]  (.A(OR4_292_Y), .B(OR4_334_Y), .C(OR4_236_Y), 
        .D(OR4_188_Y), .Y(R_DATA[1]));
    OR4 OR4_101 (.A(\R_DATA_TEMPR16[7] ), .B(\R_DATA_TEMPR17[7] ), .C(
        \R_DATA_TEMPR18[7] ), .D(\R_DATA_TEMPR19[7] ), .Y(OR4_101_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R25C0 (.BLK_EN(\BLKX0[25] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[25] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][0] ), .R_DATA({nc244, nc245, 
        \R_DATA_TEMPR25[9] , \R_DATA_TEMPR25[8] , \R_DATA_TEMPR25[7] , 
        \R_DATA_TEMPR25[6] , \R_DATA_TEMPR25[5] , \R_DATA_TEMPR25[4] , 
        \R_DATA_TEMPR25[3] , \R_DATA_TEMPR25[2] , \R_DATA_TEMPR25[1] , 
        \R_DATA_TEMPR25[0] }));
    OR4 OR4_171 (.A(\R_DATA_TEMPR24[10] ), .B(\R_DATA_TEMPR25[10] ), 
        .C(\R_DATA_TEMPR26[10] ), .D(\R_DATA_TEMPR27[10] ), .Y(
        OR4_171_Y));
    OR4 OR4_214 (.A(OR4_235_Y), .B(OR2_21_Y), .C(\R_DATA_TEMPR22[8] ), 
        .D(\R_DATA_TEMPR23[8] ), .Y(OR4_214_Y));
    OR4 OR4_246 (.A(OR4_57_Y), .B(OR4_317_Y), .C(OR4_333_Y), .D(
        OR4_31_Y), .Y(OR4_246_Y));
    OR4 OR4_221 (.A(\R_DATA_TEMPR4[3] ), .B(\R_DATA_TEMPR5[3] ), .C(
        \R_DATA_TEMPR6[3] ), .D(\R_DATA_TEMPR7[3] ), .Y(OR4_221_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R14C0 (.BLK_EN(\BLKX0[14] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[9], W_DATA[8], 
        W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], 
        W_DATA[2], W_DATA[1], W_DATA[0]}), .W_EN(\BLKZ0[14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][0] ), .R_DATA({nc246, nc247, 
        \R_DATA_TEMPR14[9] , \R_DATA_TEMPR14[8] , \R_DATA_TEMPR14[7] , 
        \R_DATA_TEMPR14[6] , \R_DATA_TEMPR14[5] , \R_DATA_TEMPR14[4] , 
        \R_DATA_TEMPR14[3] , \R_DATA_TEMPR14[2] , \R_DATA_TEMPR14[1] , 
        \R_DATA_TEMPR14[0] }));
    OR4 OR4_74 (.A(\R_DATA_TEMPR16[28] ), .B(\R_DATA_TEMPR17[28] ), .C(
        \R_DATA_TEMPR18[28] ), .D(\R_DATA_TEMPR19[28] ), .Y(OR4_74_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[1]  (.A(CFG3_0_Y), .B(CFG3_5_Y), 
        .Y(\BLKX0[1] ));
    OR4 OR4_61 (.A(OR4_165_Y), .B(OR2_19_Y), .C(\R_DATA_TEMPR22[31] ), 
        .D(\R_DATA_TEMPR23[31] ), .Y(OR4_61_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R26C2 (.BLK_EN(\BLKX0[26] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[26] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][2] ), .R_DATA({nc248, nc249, 
        \R_DATA_TEMPR26[29] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR26[27] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR26[25] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR26[23] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR26[21] , \R_DATA_TEMPR26[20] }));
    OR2 OR2_5 (.A(\R_DATA_TEMPR20[5] ), .B(\R_DATA_TEMPR21[5] ), .Y(
        OR2_5_Y));
    OR4 OR4_315 (.A(\R_DATA_TEMPR4[9] ), .B(\R_DATA_TEMPR5[9] ), .C(
        \R_DATA_TEMPR6[9] ), .D(\R_DATA_TEMPR7[9] ), .Y(OR4_315_Y));
    OR4 OR4_40 (.A(OR4_76_Y), .B(OR4_276_Y), .C(OR4_45_Y), .D(
        OR4_219_Y), .Y(OR4_40_Y));
    OR4 OR4_166 (.A(\R_DATA_TEMPR8[19] ), .B(\R_DATA_TEMPR9[19] ), .C(
        \R_DATA_TEMPR10[19] ), .D(\R_DATA_TEMPR11[19] ), .Y(OR4_166_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[28]  (.A(CFG3_21_Y), .B(
        CFG3_22_Y), .Y(\BLKX0[28] ));
    OR4 OR4_47 (.A(\R_DATA_TEMPR0[8] ), .B(\R_DATA_TEMPR1[8] ), .C(
        \R_DATA_TEMPR2[8] ), .D(\R_DATA_TEMPR3[8] ), .Y(OR4_47_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX0[23]  (.A(CFG3_15_Y), .B(
        CFG3_9_Y), .Y(\BLKX0[23] ));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R17C1 (.BLK_EN(\BLKX0[17] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][1] ), .R_DATA({nc250, nc251, 
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR17[18] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR17[16] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR17[14] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR17[12] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR17[10] }));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[3]  (.A(CFG3_23_Y), .B(CFG3_4_Y)
        , .Y(\BLKZ0[3] ));
    OR4 \OR4_R_DATA[28]  (.A(OR4_310_Y), .B(OR4_264_Y), .C(OR4_105_Y), 
        .D(OR4_143_Y), .Y(R_DATA[28]));
    OR4 OR4_98 (.A(OR4_21_Y), .B(OR2_10_Y), .C(\R_DATA_TEMPR22[23] ), 
        .D(\R_DATA_TEMPR23[23] ), .Y(OR4_98_Y));
    OR4 OR4_321 (.A(\R_DATA_TEMPR28[31] ), .B(\R_DATA_TEMPR29[31] ), 
        .C(\R_DATA_TEMPR30[31] ), .D(\R_DATA_TEMPR31[31] ), .Y(
        OR4_321_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKZ0[2]  (.A(CFG3_16_Y), .B(CFG3_4_Y)
        , .Y(\BLKZ0[2] ));
    OR4 OR4_337 (.A(OR4_46_Y), .B(OR2_35_Y), .C(\R_DATA_TEMPR22[0] ), 
        .D(\R_DATA_TEMPR23[0] ), .Y(OR4_337_Y));
    OR4 OR4_130 (.A(OR4_53_Y), .B(OR2_38_Y), .C(\R_DATA_TEMPR22[13] ), 
        .D(\R_DATA_TEMPR23[13] ), .Y(OR4_130_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R28C1 (.BLK_EN(\BLKX0[28] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[19], W_DATA[18], 
        W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], 
        W_DATA[12], W_DATA[11], W_DATA[10]}), .W_EN(\BLKZ0[28] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][1] ), .R_DATA({nc252, nc253, 
        \R_DATA_TEMPR28[19] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR28[17] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR28[15] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR28[13] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR28[11] , \R_DATA_TEMPR28[10] }));
    OR2 OR2_25 (.A(\R_DATA_TEMPR20[7] ), .B(\R_DATA_TEMPR21[7] ), .Y(
        OR2_25_Y));
    RAM64x12 LSRAM_0_PF_URAM_0_PF_URAM_R11C2 (.BLK_EN(\BLKX0[11] ), 
        .BUSY_FB(GND), .R_ADDR({R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .R_ADDR_AD_N(VCC), 
        .R_ADDR_AL_N(VCC), .R_ADDR_BYPASS(GND), .R_ADDR_EN(VCC), 
        .R_ADDR_SD(GND), .R_ADDR_SL_N(VCC), .R_CLK(CLK), .R_DATA_AD_N(
        VCC), .R_DATA_AL_N(VCC), .R_DATA_BYPASS(VCC), .R_DATA_EN(VCC), 
        .R_DATA_SD(GND), .R_DATA_SL_N(VCC), .W_ADDR({W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .W_CLK(CLK), .W_DATA({GND, GND, W_DATA[29], W_DATA[28], 
        W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], 
        W_DATA[22], W_DATA[21], W_DATA[20]}), .W_EN(\BLKZ0[11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][2] ), .R_DATA({nc254, nc255, 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR11[28] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR11[26] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR11[24] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR11[22] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR11[20] }));
    OR4 OR4_169 (.A(\R_DATA_TEMPR4[12] ), .B(\R_DATA_TEMPR5[12] ), .C(
        \R_DATA_TEMPR6[12] ), .D(\R_DATA_TEMPR7[12] ), .Y(OR4_169_Y));
    OR4 OR4_303 (.A(\R_DATA_TEMPR4[17] ), .B(\R_DATA_TEMPR5[17] ), .C(
        \R_DATA_TEMPR6[17] ), .D(\R_DATA_TEMPR7[17] ), .Y(OR4_303_Y));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
