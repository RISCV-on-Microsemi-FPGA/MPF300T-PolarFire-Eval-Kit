// Copyright 2009 Actel Corporation. All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// Revision Information:
// SVN Revision Information:
// SVN $Revision: $
module
CAHBtoAPB3OIl
(
input
wire
HCLK,
input
wire
HRESETN,
input
wire
CAHBtoAPB3Il,
input
wire
CAHBtoAPB3ll,
output
reg
PENABLE
)
;
parameter
SYNC_RESET
=
0
;
localparam
CAHBtoAPB3l0
=
2
'b
00
;
localparam
CAHBtoAPB3OOI
=
2
'b
01
;
localparam
CAHBtoAPB3IIl
=
2
'b
10
;
reg
[
1
:
0
]
CAHBtoAPB3lIl
,
CAHBtoAPB3Oll
;
reg
CAHBtoAPB3Ill
;
wire
CAHBtoAPB3O1I
;
wire
CAHBtoAPB3I1I
;
assign
CAHBtoAPB3O1I
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
HRESETN
;
assign
CAHBtoAPB3I1I
=
(
SYNC_RESET
==
1
)
?
HRESETN
:
1
'b
1
;
always
@
(
*
)
begin
CAHBtoAPB3Ill
=
1
'b
0
;
case
(
CAHBtoAPB3lIl
)
CAHBtoAPB3l0
:
begin
if
(
CAHBtoAPB3Il
)
begin
CAHBtoAPB3Oll
<=
CAHBtoAPB3OOI
;
end
else
begin
CAHBtoAPB3Oll
<=
CAHBtoAPB3l0
;
end
end
CAHBtoAPB3OOI
:
begin
CAHBtoAPB3Ill
=
1
'b
1
;
CAHBtoAPB3Oll
<=
CAHBtoAPB3IIl
;
end
CAHBtoAPB3IIl
:
begin
if
(
CAHBtoAPB3ll
)
begin
CAHBtoAPB3Oll
<=
CAHBtoAPB3l0
;
end
else
begin
CAHBtoAPB3Ill
=
1
'b
1
;
CAHBtoAPB3Oll
<=
CAHBtoAPB3IIl
;
end
end
default
:
begin
CAHBtoAPB3Ill
=
1
'b
0
;
CAHBtoAPB3Oll
<=
CAHBtoAPB3l0
;
end
endcase
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3lIl
<=
CAHBtoAPB3l0
;
PENABLE
<=
1
'b
0
;
end
else
begin
CAHBtoAPB3lIl
<=
CAHBtoAPB3Oll
;
PENABLE
<=
CAHBtoAPB3Ill
;
end
end
endmodule
