// ****************************************************************************/
// Microsemi Corporation Proprietary and Confidential
// Copyright 2015 Microsemi Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//
// Description: 
//
// SVN Revision Information:
// SVN $Revision: 25822 $
// SVN $Date: 2015-12-22 14:07:30 +0000 (Tue, 22 Dec 2015) $
//
// Resolved SARs
// SAR      Date     Who   Description
//
// Notes:
//
// ****************************************************************************/
`timescale 1ns/1ns
module testbench ();

////////////////////////////////////////////////////////////////////////////
// User modifiable parameters
////////////////////////////////////////////////////////////////////////////
parameter AXI_CLK_HALF_PERIOD = 5; // Generates an AXI CLK of 100MHz
parameter AHB_CLK_HALF_PERIOD = 5; // Generates an AHB CLK of 100MHz
parameter RAM_ADDR_WIDTH      = 7; // Determines the size of all RAM buffers
parameter RAM_INIT_FILE       = "ram_init.mem"; // MEM file containing binary
                                                // data initialise the wr_golden_mem RAM
`include "../../../../coreparameters.v"
    reg                     HCLK = 0;
    reg                     HRESETN = 0;
    wire                    HSEL;
    wire  [31:0]            HADDR;
    wire                    HWRITE;
    wire                    HREADYIN;
    wire  [1:0]             HTRANS;
    wire  [2:0]             HSIZE;
    wire  [31:0]            HWDATA;
    wire  [2:0]             HBURST;
    wire                    HMASTLOCK;
  
    wire                    HREADYOUT;
    wire                    HRESP;
    wire  [31:0]            HRDATA;
  
    reg                     ACLK = 0;
    reg                     ARESETN = 0;
    wire                    AWREADY;
    wire                    WREADY;
    wire  [ID_WIDTH-1:0]    BID;
    wire  [1:0]             BRESP;
    wire                    BVALID;
    wire                    ARREADY;
    wire  [ID_WIDTH-1:0]    RID;
    wire  [63:0]            RDATA;
    wire  [1:0]             RRESP;
    wire                    RLAST;
    wire                    RVALID;

    wire  [ID_WIDTH-1:0]    AWID;
    wire  [31:0]            AWADDR;
    wire  [3:0]             AWLEN;
    wire  [2:0]             AWSIZE;
    wire  [1:0]             AWBURST;
    wire                    AWVALID;

    wire  [ID_WIDTH-1:0]    WID;
    wire  [63:0]            WDATA;
    wire  [7:0]             WSTRB;
    wire                    WLAST;
    wire                    WVALID;
    wire                    BREADY;
    wire  [ID_WIDTH-1:0]    ARID;
    wire  [31:0]            ARADDR;
    wire  [3:0]             ARLEN;
    wire  [2:0]             ARSIZE;
    wire  [1:0]             ARBURST;
    wire                    ARVALID;
    wire                    RREADY;

// Signals normally generated by the AHB-Lite interconnect
assign HSEL = 1'b1;
assign HREADYOUT = 1'b1;
////////////////////////////////////////////////////////////////////////////////
// Clock and reset generation
////////////////////////////////////////////////////////////////////////////////
always
begin
    #AXI_CLK_HALF_PERIOD ACLK = ~ACLK;
end

always
begin
    #AHB_CLK_HALF_PERIOD HCLK = ~HCLK;
end

initial 
begin
    #100;
    HRESETN = 1'b1;
    ARESETN = 1'b1;
end

////////////////////////////////////////////////////////////////////////////////
// Instantiate DUT
////////////////////////////////////////////////////////////////////////////////
COREAXITOAHBL # (
                .ASYNC_CLOCKS       (ASYNC_CLOCKS),
                .ID_WIDTH           (ID_WIDTH),
                .NO_BURST_TRANS     (NO_BURST_TRANS),
                .WRAP_SUPPORT       (WRAP_SUPPORT)
) U_COREAXITOAHBL(
                // AXIMaster inputs
                .ACLK               (ACLK),
                .ARESETN            (ARESETN),
                .AWVALID            (AWVALID),
                .AWLEN              (AWLEN),
                .AWSIZE             (AWSIZE),
                .AWBURST            (AWBURST),
                .AWID               (AWID),
                .AWADDR             (AWADDR),
                .WVALID             (WVALID),
                .WDATA              (WDATA),
                .WSTRB              (WSTRB),
                .WLAST              (WLAST),
                .WID                (WID),
                .BREADY             (BREADY),
                .ARVALID            (ARVALID),
                .RREADY             (RREADY),
                .ARADDR             (ARADDR),
                .ARSIZE             (ARSIZE),
                .ARID               (ARID),
                .ARLEN              (ARLEN),
                .ARBURST            (ARBURST),

                // AHB Slave inputs
                .HCLK               (HCLK),
                .HRESETN            (HRESETN),
                .HREADYIN           (HREADYIN),
                .HRESP              (HRESP),
                .HRDATA             (HRDATA),

                // AXIMaster outputs
                .BRESP              (BRESP),
                .BID                (BID),
                .BVALID             (BVALID),
                .AWREADY            (AWREADY),
                .WREADY             (WREADY),
                .ARREADY            (ARREADY),
                .RVALID             (RVALID),
                .RLAST              (RLAST),
                .RID                (RID),
                .RDATA              (RDATA),
                .RRESP              (RRESP),

                // AXI Slave outputs
                .HWRITE             (HWRITE),
                .HSIZE              (HSIZE),
                .HWDATA             (HWDATA),
                .HADDR              (HADDR),
                .HTRANS             (HTRANS),
                .HBURST             (HBURST)
);   

////////////////////////////////////////////////////////////////////////////////
// Instantiate AXI Master model
////////////////////////////////////////////////////////////////////////////////
AXI_Master # (
                .ID_WIDTH           (ID_WIDTH),
                .RAM_ADDR_WIDTH     (RAM_ADDR_WIDTH),
                .RAM_INIT_FILE      (RAM_INIT_FILE)
) U_AXI_Master (
                // OUTPUT signals
                .AWREADY            (AWREADY),
                .WREADY             (WREADY),
                .BID                (BID),
                .BRESP              (BRESP),
                .BVALID             (BVALID),
                .ARREADY            (ARREADY),
                .RID                (RID),
                .RDATA              (RDATA),
                .RRESP              (RRESP),
                .RLAST              (RLAST),
                .RVALID             (RVALID),

                // INPUT signals
                .ACLK               (ACLK),
                .ARESETN            (ARESETN),
                .AWID               (AWID),
                .AWADDR             (AWADDR),
                .AWLEN              (AWLEN),
                .AWSIZE             (AWSIZE),
                .AWBURST            (AWBURST),
                .AWVALID            (AWVALID),
                .WID                (WID),
                .WDATA              (WDATA),
                .WSTRB              (WSTRB),
                .WLAST              (WLAST),
                .WVALID             (WVALID),
                .BREADY             (BREADY),
                .ARID               (ARID),
                .ARADDR             (ARADDR),
                .ARLEN              (ARLEN),
                .ARSIZE             (ARSIZE),
                .ARBURST            (ARBURST),
                .ARVALID            (ARVALID),
                .RREADY             (RREADY)
);

////////////////////////////////////////////////////////////////////////////////
// Instantiate AHB Slave BFM
////////////////////////////////////////////////////////////////////////////////
AHBL_Slave # (
                .RAM_ADDR_WIDTH     (RAM_ADDR_WIDTH)
) U_AHBL_Slave (
                .HCLK               (HCLK),
                .HRESETN            (HRESETN),
                .HWRITE             (HWRITE),
                .HSEL               (HSEL),
                .HTRANS             (HTRANS),
                .HSIZE              (HSIZE),
                .HADDR              (HADDR),
                .HBURST             (HBURST),
                .HWDATA             (HWDATA),
                .HMASTLOCK          (HMASTLOCK), 
                .HREADY_slave       (HREADYOUT),

                .HREADYOUT_slave    (HREADYIN),
                .HRESP              (HRESP),
                .HRDATA             (HRDATA)
);

endmodule // testbench
