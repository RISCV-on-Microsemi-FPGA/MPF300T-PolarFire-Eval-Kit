// Copyright 2009 Actel Corporation. All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// Revision Information:
// SVN Revision Information:
// SVN $Revision: $
module
COREAHBTOAPB3
(
input
wire
HCLK,
input
wire
HRESETN,
input
wire
HSEL,
input
wire
[
31
:
0
]
HADDR,
input
wire
HWRITE,
input
wire
HREADY,
input
wire
[
1
:
0
]
HTRANS,
input
wire
[
31
:
0
]
HWDATA,
output
wire
HREADYOUT,
output
wire
[
1
:
0
]
HRESP,
output
wire
[
31
:
0
]
HRDATA,
output
wire
[
31
:
0
]
PADDR,
output
wire
PWRITE,
output
wire
PENABLE,
output
wire
[
31
:
0
]
PWDATA,
output
wire
PSEL,
input
wire
PREADY,
input
wire
PSLVERR,
input
wire
[
31
:
0
]
PRDATA
)
;
parameter
FAMILY
=
17
;
parameter
SYNC_RESET
=
(
FAMILY
==
25
)
?
1
:
0
;
wire
CAHBtoAPB3Il
;
wire
CAHBtoAPB3ll
;
wire
CAHBtoAPB3l
;
wire
CAHBtoAPB3OI
;
wire
CAHBtoAPB3II
;
wire
CAHBtoAPB3lI
;
wire
CAHBtoAPB3Ol
;
CAHBtoAPB3O
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBtoAPB3lll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.HSEL
(
HSEL
)
,
.CAHBtoAPB3I
(
HTRANS
[
1
]
)
,
.HWRITE
(
HWRITE
)
,
.HREADY
(
HREADY
)
,
.HRESP
(
HRESP
)
,
.HREADYOUT
(
HREADYOUT
)
,
.PREADY
(
PREADY
)
,
.PSLVERR
(
PSLVERR
)
,
.PENABLE
(
PENABLE
)
,
.PWRITE
(
PWRITE
)
,
.PSEL
(
PSEL
)
,
.CAHBtoAPB3l
(
CAHBtoAPB3l
)
,
.CAHBtoAPB3OI
(
CAHBtoAPB3OI
)
,
.CAHBtoAPB3II
(
CAHBtoAPB3II
)
,
.CAHBtoAPB3lI
(
CAHBtoAPB3lI
)
,
.CAHBtoAPB3Ol
(
CAHBtoAPB3Ol
)
,
.CAHBtoAPB3Il
(
CAHBtoAPB3Il
)
,
.CAHBtoAPB3ll
(
CAHBtoAPB3ll
)
)
;
CAHBtoAPB3OIl
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBtoAPB3O0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBtoAPB3Il
(
CAHBtoAPB3Il
)
,
.CAHBtoAPB3ll
(
CAHBtoAPB3ll
)
,
.PENABLE
(
PENABLE
)
)
;
CAHBtoAPB3l1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBtoAPB3I0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBtoAPB3l
(
CAHBtoAPB3l
)
,
.CAHBtoAPB3OI
(
CAHBtoAPB3OI
)
,
.CAHBtoAPB3II
(
CAHBtoAPB3II
)
,
.CAHBtoAPB3lI
(
CAHBtoAPB3lI
)
,
.CAHBtoAPB3Ol
(
CAHBtoAPB3Ol
)
,
.HADDR
(
HADDR
[
31
:
0
]
)
,
.HWDATA
(
HWDATA
[
31
:
0
]
)
,
.HRDATA
(
HRDATA
[
31
:
0
]
)
,
.PADDR
(
PADDR
[
31
:
0
]
)
,
.PWDATA
(
PWDATA
[
31
:
0
]
)
,
.PRDATA
(
PRDATA
[
31
:
0
]
)
)
;
endmodule
