// Copyright 2009 Actel Corporation. All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// Revision Information:
// SVN Revision Information:
// SVN $Revision: $
module
CAHBtoAPB3l1I
(
input
wire
HCLK,
input
wire
HRESETN,
input
wire
CAHBtoAPB3l,
input
wire
CAHBtoAPB3OI,
input
wire
CAHBtoAPB3II,
input
wire
CAHBtoAPB3lI,
input
wire
CAHBtoAPB3Ol,
input
wire
[
31
:
0
]
HADDR,
input
wire
[
31
:
0
]
HWDATA,
output
reg
[
31
:
0
]
HRDATA,
output
reg
[
31
:
0
]
PADDR,
output
reg
[
31
:
0
]
PWDATA,
input
wire
[
31
:
0
]
PRDATA
)
;
parameter
SYNC_RESET
=
0
;
reg
[
31
:
0
]
CAHBtoAPB3OOl
;
reg
[
31
:
0
]
CAHBtoAPB3IOl
;
reg
[
31
:
0
]
CAHBtoAPB3lOl
;
wire
CAHBtoAPB3O1I
;
wire
CAHBtoAPB3I1I
;
assign
CAHBtoAPB3O1I
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
HRESETN
;
assign
CAHBtoAPB3I1I
=
(
SYNC_RESET
==
1
)
?
HRESETN
:
1
'b
1
;
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3OOl
<=
32
'b
0
;
end
else
begin
if
(
CAHBtoAPB3l
)
begin
CAHBtoAPB3OOl
<=
HADDR
[
31
:
0
]
;
end
else
begin
if
(
CAHBtoAPB3Ol
)
begin
CAHBtoAPB3OOl
<=
CAHBtoAPB3IOl
[
31
:
0
]
;
end
end
end
end
always
@
(
*
)
begin
PADDR
=
CAHBtoAPB3OOl
[
31
:
0
]
;
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3IOl
<=
32
'b
0
;
end
else
begin
if
(
CAHBtoAPB3lI
)
begin
CAHBtoAPB3IOl
<=
HADDR
[
31
:
0
]
;
end
end
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
CAHBtoAPB3lOl
<=
32
'b
0
;
end
else
begin
if
(
CAHBtoAPB3OI
)
begin
CAHBtoAPB3lOl
[
31
:
0
]
<=
HWDATA
[
31
:
0
]
;
end
end
end
always
@
(
*
)
begin
PWDATA
[
31
:
0
]
=
CAHBtoAPB3lOl
[
31
:
0
]
;
end
always
@
(
posedge
HCLK
or
negedge
CAHBtoAPB3O1I
)
begin
if
(
(
!
CAHBtoAPB3O1I
)
||
(
!
CAHBtoAPB3I1I
)
)
begin
HRDATA
[
31
:
0
]
<=
32
'b
0
;
end
else
begin
if
(
CAHBtoAPB3II
)
begin
HRDATA
[
31
:
0
]
<=
PRDATA
[
31
:
0
]
;
end
end
end
endmodule
